{"andra|NUM": 1000000.0, "arton|NUM": 1000000.0, "bakre|ADJ": 1000000.0, "brunch|NOUN": 1000000.0, "decimeter|NOUN": 1000000.0, "elva|NUM": 1000000.0, "ett|NUM": 1000000.0, "Europa|PROPN": 1000000.0, "fem|NUM": 1000000.0, "femte|NUM": 1000000.0, "femtio|NUM": 1000000.0, "femton|NUM": 1000000.0, "fjorton|NUM": 1000000.0, "fjärde|NUM": 1000000.0, "främre|ADJ": 1000000.0, "fyra|NUM": 1000000.0, "fyrtio|NUM": 1000000.0, "första|NUM": 1000000.0, "Grekland|PROPN": 1000000.0, "Göteborg|PROPN": 1000000.0, "hekto|NOUN": 1000000.0, "hela|NOUN": 1000000.0, "hundra|NUM": 1000000.0, "hundratusen|NUM": 1000000.0, "hörsel|NOUN": 1000000.0, "inrikesminister|NOUN": 1000000.0, "inrikespolitik|NOUN": 1000000.0, "Italien|PROPN": 1000000.0, "Kina|PROPN": 1000000.0, "kvällsmål|NOUN": 1000000.0, "känsel|NOUN": 1000000.0, "mellanmål|NOUN": 1000000.0, "miljard|NUM": 1000000.0, "miljon|NUM": 1000000.0, "milligram|NOUN": 1000000.0, "millimeter|NOUN": 1000000.0, "morbror|NOUN": 1000000.0, "månadsskifte|NOUN": 1000000.0, "nia|NOUN": 1000000.0, "nio|NUM": 1000000.0, "nionde|NUM": 1000000.0, "nittio|NUM": 1000000.0, "nitton|NUM": 1000000.0, "nordost|NOUN": 1000000.0, "Norge|PROPN": 1000000.0, "pingst|NOUN": 1000000.0, "Polen|PROPN": 1000000.0, "Ryssland|PROPN": 1000000.0, "sex|NUM": 1000000.0, "sexa|NOUN": 1000000.0, "sextio|NUM": 1000000.0, "sexton|NUM": 1000000.0, "sju|NUM": 1000000.0, "sjua|NOUN": 1000000.0, "sjunde|NUM": 1000000.0, "sjuttio|NUM": 1000000.0, "sjutton|NUM": 1000000.0, "sjätte|NUM": 1000000.0, "Stockholm|PROPN": 1000000.0, "storasyster|NOUN": 1000000.0, "Storbritannien|PROPN": 1000000.0, "syd|NOUN": 1000000.0, "sydväst|NOUN": 1000000.0, "sydöst|NOUN": 1000000.0, "syssling|NOUN": 1000000.0, "tia|NOUN": 1000000.0, "tio|NUM": 1000000.0, "tionde|NUM": 1000000.0, "tiotusen|NUM": 1000000.0, "tjugo|NUM": 1000000.0, "tolv|NUM": 1000000.0, "tre|NUM": 1000000.0, "tredje|NUM": 1000000.0, "trettio|NUM": 1000000.0, "tretton|NUM": 1000000.0, "tusen|NUM": 1000000.0, "två|NUM": 1000000.0, "utbildningsminister|NOUN": 1000000.0, "veckodag|NOUN": 1000000.0, "åtta|NOUN": 1000000.0, "åtta|NUM": 1000000.0, "åttio|NUM": 1000000.0, "åttonde|NUM": 1000000.0, "änkeman|NOUN": 1000000.0, "änkling|NOUN": 1000000.0, "ögonlock|NOUN": 1000000.0, "och (vardagl. å; förk. o.)|CCONJ": 26019.68, "vara (vardagl. va)|VERB": 23017.26, "i|ADP": 19272.89, "ha|VERB": 15983.31, "dess|PRON": 15935.58, "det|PRON": 14582.21, "en|DET": 14511.22, "som|PRON": 12734.7, "på|ADP": 12591.15, "å|ADP": 12462.73, "av|ADP": 11540.13, "för|ADP": 11408.82, "att|SCONJ": 11271.57, "kunna|VERB": 11119.08, "skola|AUX": 10411.19, "jag|PRON": 9390.67, "inte (formellt: icke, ej)|ADV": 9073.55, "med|ADP": 8790.85, "till|ADP": 8662.68, "liten|ADJ": 8654.67, "den|DET": 6896.18, "ett|DET": 6314.26, "analog|ADJ": 5649.0, "unna|VERB": 5559.15, "om|ADP": 5278.24, "vi|PRON": 4723.57, "men|CCONJ": 4545.97, "man|PRON": 4446.34, "de (vardagl. dom)|DET": 4437.26, "få|VERB": 4060.39, "så|ADV": 4004.97, "som|CCONJ": 3762.28, "sig (vardagl. sej)|PRON": 3469.03, "han|PRON": 3380.88, "de (vardagl. dom)|PRON": 3345.8, "bli|VERB": 3293.35, "komma|VERB": 3224.74, "det|DET": 3221.41, "sin|PRON": 3217.3, "eller|CCONJ": 3138.92, "från|ADP": 3117.46, "mycket|ADV": 3112.13, "vilja|VERB": 3004.91, "all|PRON": 2975.47, "göra|VERB": 2942.04, "om|SCONJ": 2630.45, "annan|PRON": 2624.2, "du|PRON": 2581.46, "någon (vardagl. nån, förk. ngn)|PRON": 2565.69, "finna|VERB": 2465.41, "ta (el. taga)|VERB": 2452.4, "när|ADV": 2386.89, "se|VERB": 2253.32, "måste|AUX": 2214.95, "detta|PRON": 2200.74, "stor|ADJ": 2046.73, "nu|ADV": 2033.06, "gå|VERB": 2001.14, "säga|VERB": 1998.46, "den|PRON": 1981.49, "vad (vardagl. va)|PRON": 1911.2, "år|NOUN": 1886.72, "äga|VERB": 1867.88, "under|ADP": 1851.63, "betyda|VERB": 1811.72, "också (vardagl. oxå)|ADV": 1797.39, "där|ADV": 1790.68, "då|ADV": 1788.93, "min|PRON": 1757.18, "böra|AUX": 1743.31, "hur|ADV": 1690.32, "mig (vardagl. mej)|PRON": 1622.7, "mot|ADP": 1592.42, "bara|ADV": 1582.15, "vilken|PRON": 1512.84, "ut|ADV": 1481.5, "ny|ADJ": 1446.08, "vid|ADP": 1439.02, "än|CCONJ": 1428.89, "bra|ADJ": 1428.27, "ingen|PRON": 1350.9, "dem (vardagl. dom)|PRON": 1341.39, "efter|ADP": 1323.97, "upp|PART": 1322.38, "hon|PRON": 1291.75, "lite|ADV": 1288.09, "denna|PRON": 1279.97, "in|ADV": 1274.61, "mycket|ADJ": 1271.67, "över|ADP": 1267.18, "ge (formellt giva)|VERB": 1208.51, "vår (vardagl. våran)|PRON": 1206.78, "del|NOUN": 1202.45, "här|ADV": 1194.91, "även|ADV": 1191.77, "skriva|VERB": 1141.32, "tid|NOUN": 1127.59, "ju|ADV": 1119.58, "sedan (vardagl. sen)|ADV": 1115.12, "te sig|VERB": 1115.09, "riva|VERB": 1088.02, "börja|VERB": 1039.45, "hel|ADJ": 1034.76, "dag|NOUN": 1033.61, "själv|PRON": 1033.19, "människa|NOUN": 1030.33, "land|NOUN": 949.12, "svensk|ADJ": 948.52, "fråga|NOUN": 938.78, "oss|PRON": 934.32, "tro|VERB": 928.39, "el|NOUN": 925.85, "tycka|VERB": 924.85, "kommentar|NOUN": 924.68, "veta|VERB": 894.31, "idag (el. i dag)|ADV": 865.13, "försöka|VERB": 859.72, "behöva|VERB": 858.16, "samma|PRON": 844.13, "mellan|ADP": 841.51, "känna|VERB": 840.25, "läsa|VERB": 823.05, "ro|VERB": 816.02, "kanske|ADV": 809.75, "lik|ADJ": 808.09, "låta|VERB": 807.17, "olik|ADJ": 790.47, "sådan|PRON": 788.97, "sätt|NOUN": 784.91, "hans|PRON": 774.6, "din|PRON": 771.62, "gång|NOUN": 763.39, "stå|VERB": 761.8, "inom|ADP": 758.15, "visa|VERB": 757.44, "använda|VERB": 749.26, "vända|VERB": 749.26, "hålla|VERB": 739.42, "genom|ADP": 733.74, "helt|ADV": 721.67, "fler|ADJ": 717.99, "utan|ADP": 707.53, "väl|ADV": 705.75, "barn|NOUN": 700.31, "enligt|ADP": 680.22, "tänka|VERB": 666.7, "ni|PRON": 665.01, "viktig|ADJ": 662.11, "ring|NOUN": 658.84, "eftersom|SCONJ": 652.0, "liv|NOUN": 624.66, "deras|PRON": 623.86, "värld|NOUN": 617.89, "viss|ADJ": 614.61, "dock|ADV": 614.54, "egen|ADJ": 612.48, "folk|NOUN": 606.98, "regering|NOUN": 603.37, "fram|PART": 600.53, "honom|PRON": 597.56, "söka|VERB": 596.07, "dig (vardagl. dej)|PRON": 590.81, "utan|CCONJ": 586.71, "sak|NOUN": 581.51, "hög|ADJ": 578.03, "länge|ADV": 568.83, "person|NOUN": 568.43, "ligga|VERB": 566.6, "son|NOUN": 560.93, "både|CCONJ": 554.95, "just|ADV": 545.57, "lägga|VERB": 545.17, "antal|NOUN": 542.86, "redan|ADV": 533.67, "kvinna|NOUN": 521.11, "problem|NOUN": 520.62, "fall|NOUN": 520.07, "man|NOUN": 520.07, "aldrig|ADV": 511.81, "ofta|ADV": 501.79, "varje|DET": 501.7, "artikel|NOUN": 501.28, "anse|VERB": 500.58, "öva|VERB": 496.12, "lag|NOUN": 380.83, "slag|NOUN": 487.59, "tal|NOUN": 485.93, "åt|ADP": 484.56, "nog|ADV": 482.6, "bok|NOUN": 478.59, "varför|ADV": 475.84, "handla|VERB": 475.07, "gammal|ADJ": 470.38, "bild|NOUN": 468.8, "sida|NOUN": 466.09, "så|SCONJ": 465.43, "öka|VERB": 462.83, "därför|ADV": 461.58, "sen|ADJ": 459.09, "god|ADJ": 453.87, "hos|ADP": 453.15, "alltid|ADV": 446.85, "skapa|VERB": 445.51, "arbete|NOUN": 441.9, "kapa|VERB": 435.8, "samt|CCONJ": 435.23, "blogg|NOUN": 430.91, "innan|SCONJ": 429.65, "som|ADV": 429.24, "ur|ADP": 427.0, "gälla|VERB": 426.9, "verka|VERB": 423.62, "tala|VERB": 423.1, "bära|VERB": 422.35, "för|ADV": 421.08, "väg|NOUN": 420.51, "samhälle|NOUN": 420.38, "alltså|ADV": 419.06, "stat|NOUN": 416.16, "stad|NOUN": 413.66, "höra|VERB": 412.78, "innebära|VERB": 412.65, "genom att|SCONJ": 412.39, "företag|NOUN": 412.18, "möjlighet|NOUN": 411.21, "ord|NOUN": 410.3, "politisk|ADJ": 409.23, "välja|VERB": 403.72, "er|PRON": 403.6, "förstå|VERB": 403.12, "inlägg|NOUN": 403.03, "ägg|NOUN": 403.03, "te|NOUN": 401.97, "spela|VERB": 401.87, "så att|SCONJ": 400.31, "lika|ADV": 394.25, "hitta|VERB": 390.73, "tag|NOUN": 390.12, "dra|VERB": 389.89, "leda|VERB": 388.53, "gärna|ADV": 387.27, "ändå|ADV": 386.11, "förslag|NOUN": 385.31, "lyckas|VERB": 384.14, "dessutom|ADV": 381.45, "område|NOUN": 380.95, "svår|ADJ": 379.67, "lära|VERB": 376.66, "sätta|VERB": 375.3, "plats|NOUN": 374.33, "lång|ADJ": 372.0, "lämna|VERB": 369.7, "bygga|VERB": 368.34, "politik|NOUN": 367.14, "tidigare|ADV": 366.98, "kalla|VERB": 365.74, "peng|NOUN": 365.1, "väldigt|ADV": 363.6, "leva|VERB": 363.55, "ställa|VERB": 361.06, "följa|VERB": 359.7, "vecka|NOUN": 357.71, "ja|INTJ": 353.15, "ske|VERB": 351.8, "parti|NOUN": 348.11, "kräva|VERB": 347.5, "utveckling|NOUN": 341.81, "faktiskt|ADV": 341.44, "ena|VERB": 340.46, "svara|VERB": 339.8, "ner|PART": 339.66, "fortsätta|VERB": 337.29, "skola|NOUN": 334.72, "bruka|VERB": 334.18, "mål|NOUN": 331.84, "par|NOUN": 331.61, "sent|ADV": 330.39, "ekonomisk|ADJ": 327.88, "kl. (klockan)|NOUN": 325.82, "dålig|ADJ": 323.94, "namn|NOUN": 323.21, "igen|ADV": 321.76, "verkligen|ADV": 321.76, "mena|VERB": 320.45, "fortfarande|ADV": 319.39, "grupp|NOUN": 315.91, "beslut|NOUN": 315.74, "även om|SCONJ": 314.71, "enda|ADJ": 314.53, "bort|PART": 313.64, "slå|VERB": 312.71, "möjlig|ADJ": 310.72, "många|PRON": 310.01, "hända|VERB": 307.66, "ämna|AUX": 307.66, "endast|ADV": 302.17, "miljon|NOUN": 301.59, "vidare|ADV": 297.7, "ganska|ADV": 295.35, "svar|NOUN": 291.65, "varenda|DET": 291.39, "istället (el. i stället)|ADV": 291.38, "först|ADV": 290.35, "arbeta|VERB": 289.93, "heller|ADV": 288.81, "riktigt|ADV": 288.62, "hand|NOUN": 288.6, "uppgift|NOUN": 287.98, "fungera (vardagl. funka)|VERB": 287.4, "beta|VERB": 286.58, "köpa|VERB": 284.11, "nästan|ADV": 284.0, "bra|ADV": 283.65, "bland|ADP": 282.47, "december|NOUN": 280.83, "sitta|VERB": 280.32, "precis|ADV": 277.18, "hennes|PRON": 275.94, "åta sig|VERB": 275.39, "bland annat (förk. bl.a.)|ADV": 275.2, "krig|NOUN": 275.09, "till exempel (förk. t.ex., t ex)|ADV": 274.97, "tillsammans|ADV": 274.88, "henne|PRON": 272.82, "intressant|ADJ": 272.16, "val|NOUN": 13.73, "kyrka|NOUN": 268.45, "egentligen|ADV": 267.44, "inför|ADP": 267.33, "historia|NOUN": 267.25, "jobb|NOUN": 266.97, "berätta|VERB": 266.34, "vanlig|ADJ": 265.84, "rätta|VERB": 265.36, "januari|NOUN": 264.41, "information|NOUN": 264.14, "flest|ADJ": 262.77, "ung|ADJ": 260.53, "en|PRON": 260.31, "tillbaka (vardagl. tillbaks)|PART": 259.58, "film|NOUN": 258.67, "ibland (el. i bland)|ADV": 258.58, "medan (vardagl. medans)|SCONJ": 257.43, "slut|NOUN": 256.6, "massa|NOUN": 255.87, "tanke|NOUN": 251.61, "akt|NOUN": 251.45, "procent|NOUN": 251.21, "månad|NOUN": 251.14, "sista|ADJ": 250.04, "ätt|NOUN": 249.91, "sluta|VERB": 249.47, "verksamhet|NOUN": 249.2, "rätt|NOUN": 249.15, "samtidigt|ADV": 247.54, "emot|ADP": 247.28, "stöd|NOUN": 244.26, "familj|NOUN": 244.19, "vem|PRON": 243.27, "åka|VERB": 243.14, "betala|VERB": 242.04, "kommun|NOUN": 242.01, "resultat|NOUN": 241.96, "utveckla|VERB": 241.91, "föra|VERB": 240.44, "hjälpa|VERB": 238.92, "nästa|ADJ": 237.94, "nära|ADV": 237.62, "nej|INTJ": 237.61, "text|NOUN": 234.6, "exempel|NOUN": 232.43, "särskilt|ADV": 232.35, "debatt|NOUN": 232.07, "när det gäller|ADP": 230.03, "på grund av (förk. p.g.a, pga., p g a)|ADV": 229.03, "situation|NOUN": 229.02, "europeisk|ADJ": 228.56, "form|NOUN": 228.11, "orm|NOUN": 228.11, "råd|NOUN": 228.07, "november|NOUN": 228.05, "makt|NOUN": 228.02, "social|ADJ": 226.91, "vinna|VERB": 226.63, "kvar|PART": 226.35, "system|NOUN": 225.72, "vänta|VERB": 225.55, "tidig|ADJ": 225.46, "åtgärd|NOUN": 223.86, "krav|NOUN": 223.66, "skillnad|NOUN": 223.65, "riksdag|NOUN": 223.14, "internationell|ADJ": 222.66, "nationell|ADJ": 222.66, "jobba|VERB": 221.99, "klara|VERB": 218.16, "typ|NOUN": 217.75, "kring|ADP": 217.05, "båda (vardagl. bägge)|PRON": 217.0, "cirka (förk. ca)|ADV": 216.97, "tur|NOUN": 216.52, "polis|NOUN": 216.42, "medium|NOUN": 215.79, "låg|ADJ": 214.24, "varandra (vardagl. varann)|PRON": 214.16, "mun|NOUN": 213.93, "ansvar|NOUN": 213.48, "roll|NOUN": 213.39, "regel|NOUN": 211.92, "oktober|NOUN": 211.56, "prata|VERB": 211.06, "organisation|NOUN": 210.61, "medlem|NOUN": 210.54, "fråga|VERB": 210.47, "anmäla|VERB": 209.8, "nå|VERB": 209.69, "bo|VERB": 209.48, "krona|NOUN": 207.79, "stämma|VERB": 207.42, "rättighet|NOUN": 207.42, "sedan (vardagl. sen)|ADP": 207.3, "bakom|ADP": 206.72, "efter att|SCONJ": 206.69, "därmed|ADV": 206.58, "med|ADV": 206.58, "hus|NOUN": 206.57, "vän|NOUN": 205.79, "dela|VERB": 205.43, "februari|NOUN": 205.04, "kort|ADJ": 204.59, "grund|NOUN": 204.34, "runt|ADP": 203.5, "framtid|NOUN": 203.16, "köra|VERB": 203.16, "etikett|NOUN": 202.31, "fri|ADJ": 201.84, "behov|NOUN": 201.71, "timme (el. timma)|NOUN": 201.49, "september|NOUN": 201.31, "hoppas|VERB": 200.99, "ensam|ADJ": 200.63, "snart|ADV": 199.9, "rätt|ADV": 198.64, "förklara|VERB": 198.04, "ledning|NOUN": 197.93, "intresse|NOUN": 197.41, "tvinga|VERB": 196.99, "påverka|VERB": 196.4, "anledning|NOUN": 195.88, "titta|VERB": 195.79, "minska|VERB": 195.42, "i alla fall (el. iallafall; förk. iaf)|ADV": 195.28, "däremot|ADV": 194.9, "direkt|ADV": 194.63, "ekonomi|NOUN": 194.28, "bestämma|VERB": 192.88, "skicka|VERB": 192.84, "trots|ADP": 192.43, "åsikt|NOUN": 192.3, "diskussion|NOUN": 192.14, "rad|NOUN": 192.14, "faktum|NOUN": 192.11, "tidning|NOUN": 191.91, "mening|NOUN": 191.16, "utanför|ADP": 190.63, "rätt|ADJ": 190.49, "gemensam|ADJ": 189.45, "klar|ADJ": 187.9, "juni|NOUN": 186.95, "is|NOUN": 186.84, "bil|NOUN": 186.44, "myndighet|NOUN": 186.22, "nummer (förk. nr)|NOUN": 186.0, "allmän|ADJ": 185.28, "musik|NOUN": 185.07, "ändra|VERB": 184.81, "träffa|VERB": 184.74, "ihop|PART": 183.73, "diskutera|VERB": 183.54, "driva|VERB": 183.3, "sälja|VERB": 182.71, "sakna|VERB": 182.57, "program|NOUN": 182.39, "ifrån|ADP": 181.44, "länka|VERB": 179.35, "kunskap|NOUN": 179.19, "snabbt|ADV": 178.68, "maj|NOUN": 177.76, "amerikansk|ADJ": 177.66, "tyda|VERB": 177.46, "särskild|ADJ": 177.43, "början|NOUN": 176.59, "naturligtvis|ADV": 176.31, "skäl|NOUN": 175.99, "fin|ADJ": 174.99, "genomföra|VERB": 174.86, "liksom|ADV": 174.75, "via|ADP": 174.12, "före|ADP": 173.85, "dom|NOUN": 173.6, "risk|NOUN": 173.27, "enkel|ADJ": 173.1, "alls|ADV": 173.06, "pris|NOUN": 172.92, "räkna|VERB": 172.91, "beskriva|VERB": 172.36, "hem|PART": 172.22, "möta|VERB": 172.02, "såsom|SCONJ": 171.86, "idé|NOUN": 171.57, "gram|NOUN": 171.53, "förra|ADJ": 170.92, "tjänst|NOUN": 170.63, "heta|VERB": 170.22, "kultur|NOUN": 170.1, "äta|VERB": 169.74, "syfte|NOUN": 168.82, "princip|NOUN": 167.86, "flytta|VERB": 167.68, "ute|ADV": 167.61, "utgöra|VERB": 167.61, "politiker|NOUN": 167.43, "lätt|ADJ": 167.41, "förälder|NOUN": 167.0, "marknad|NOUN": 166.13, "nämligen|ADV": 165.98, "tydlig|ADJ": 165.93, "utbildning|NOUN": 165.87, "röra|VERB": 165.68, "nivå|NOUN": 165.64, "april|NOUN": 165.36, "mängd|NOUN": 165.27, "betydelse|NOUN": 165.2, "kristen|ADJ": 164.51, "dö|VERB": 164.3, "mars|NOUN": 164.22, "allt|ADV": 163.95, "kväll|NOUN": 163.87, "bildning|NOUN": 163.82, "länk|NOUN": 163.54, "växa|VERB": 162.65, "per|ADP": 162.15, "offentlig|ADJ": 161.83, "såväl|CCONJ": 161.72, "våga|VERB": 161.66, "vatten|NOUN": 161.3, "håll|NOUN": 161.22, "mänsklig|ADJ": 160.58, "demokrati|NOUN": 160.56, "fatta|VERB": 160.43, "jord|NOUN": 159.88, "känsla|NOUN": 159.45, "förändring|NOUN": 159.43, "nämna|VERB": 159.17, "tyvärr|ADV": 159.15, "enskild|ADJ": 159.02, "rätt|PART": 158.98, "be (el. bedja)|VERB": 158.82, "punkt|NOUN": 158.58, "ändring|NOUN": 158.58, "mission|NOUN": 158.08, "igår (el. i går)|ADV": 157.53, "kommission|NOUN": 157.33, "ort|NOUN": 156.85, "anta|VERB": 156.58, "trots att|SCONJ": 156.41, "spel|NOUN": 156.33, "språk|NOUN": 156.31, "föreslå|VERB": 156.27, "igenom|ADP": 154.93, "undra|VERB": 154.38, "eget|ADJ": 154.19, "möte|NOUN": 153.97, "mat|NOUN": 153.94, "gräns|NOUN": 153.55, "lyssna|VERB": 152.94, "delta|VERB": 152.8, "samarbete|NOUN": 152.7, "annars|ADV": 152.6, "falla|VERB": 152.58, "nära|ADJ": 152.36, "rum|NOUN": 152.07, "ungefär|ADV": 151.93, "starta|VERB": 151.68, "inse|VERB": 151.51, "internet|NOUN": 151.38, "hov|NOUN": 150.99, "öppen|ADJ": 150.86, "bidra|VERB": 150.84, "död|NOUN": 150.59, "luta|VERB": 150.2, "öga|NOUN": 150.07, "säkert|ADV": 149.46, "ämne|NOUN": 149.25, "få|ADJ": 148.91, "augusti|NOUN": 148.76, "socialdemokrat (vardagl. sosse)|NOUN": 148.49, "projekt|NOUN": 148.31, "övrig|ADJ": 148.21, "dels|CCONJ": 148.09, "framför allt (el. framförallt)|ADV": 147.43, "positiv|ADJ": 147.36, "rolig|ADJ": 147.33, "port|NOUN": 146.95, "bero|VERB": 146.68, "kropp|NOUN": 145.82, "minnas|VERB": 145.43, "handling|NOUN": 145.37, "rösta|VERB": 145.06, "riktig|ADJ": 144.98, "rapport|NOUN": 144.86, "lösning|NOUN": 144.58, "personlig|ADJ": 143.81, "kommentera|VERB": 142.95, "som att|SCONJ": 142.78, "gilla|VERB": 142.42, "bryta|VERB": 142.11, "hjälp|NOUN": 142.06, "juli|NOUN": 142.01, "innehålla|VERB": 141.45, "liknande|ADJ": 140.93, "tillfälle|NOUN": 140.9, "inte ens|ADV": 140.79, "känd|ADJ": 140.65, "forskning|NOUN": 140.49, "kraft|NOUN": 140.46, "helt enkelt|ADV": 140.11, "brott|NOUN": 139.94, "exempelvis|ADV": 139.94, "röst|NOUN": 139.89, "bjuda|VERB": 139.86, "till och med (förk. t.o.m., t o m)|ADV": 139.7, "hävda|VERB": 139.57, "hamna|VERB": 139.4, "effekt|NOUN": 138.78, "enhet|NOUN": 138.39, "det vill säga (förk. d.v.s., dvs.)|ADV": 138.07, "kontakt|NOUN": 137.86, "takt|NOUN": 137.86, "värde|NOUN": 137.82, "förutsättning|NOUN": 137.72, "sats|NOUN": 137.65, "medlemsstat|NOUN": 137.58, "hinna|VERB": 137.35, "sanning|NOUN": 136.75, "religion|NOUN": 136.55, "källa|NOUN": 136.13, "må|VERB": 135.98, "kostnad|NOUN": 135.72, "medborgare|NOUN": 135.65, "förhållande|NOUN": 135.64, "far (el. fader, vardagl. farsa)|NOUN": 135.06, "miljard|NOUN": 134.96, "ungdom|NOUN": 134.37, "släppa|VERB": 134.32, "enbart|ADV": 134.15, "drag|NOUN": 134.15, "verklighet|NOUN": 133.94, "författare|NOUN": 133.87, "tillgång|NOUN": 133.5, "nödvändig|ADJ": 133.42, "full|ADJ": 133.12, "frihet|NOUN": 132.47, "passa|VERB": 132.39, "lokal|ADJ": 132.16, "ytterligare|ADV": 131.58, "öppna|VERB": 131.53, "införa|VERB": 130.26, "ledare|NOUN": 129.98, "mamma|NOUN": 129.87, "sammanhang|NOUN": 129.67, "svensk|NOUN": 129.62, "hemma|ADV": 129.59, "produkt|NOUN": 129.58, "därefter|ADV": 129.33, "efter|ADV": 129.33, "match|NOUN": 129.11, "tro|NOUN": 129.11, "alldeles|ADV": 128.37, "lätt|ADV": 128.34, "sann|ADJ": 128.33, "uppfattning|NOUN": 128.3, "demokrat|NOUN": 128.13, "bolag|NOUN": 128.01, "erfarenhet|NOUN": 127.97, "kritik|NOUN": 127.81, "grad|NOUN": 127.76, "jude|NOUN": 127.57, "vacker|ADJ": 127.57, "erbjuda|VERB": 127.44, "kamp|NOUN": 127.43, "period|NOUN": 127.37, "modern|ADJ": 127.04, "spelare|NOUN": 127.02, "elev|NOUN": 127.01, "utredning|NOUN": 126.93, "ingå|VERB": 126.92, "kung|NOUN": 126.7, "bestå|VERB": 126.46, "katt|NOUN": 126.45, "konstatera|VERB": 126.41, "dit|ADV": 126.29, "klart|ADV": 126.22, "nuvarande|ADJ": 126.21, "styra|VERB": 126.2, "förlora|VERB": 126.19, "vit|ADJ": 126.15, "klocka|NOUN": 125.96, "påstå|VERB": 125.75, "skatt|NOUN": 125.65, "besluta|VERB": 125.13, "befolkning|NOUN": 125.01, "avse|VERB": 124.91, "ro|NOUN": 124.53, "privat|ADJ": 124.48, "steg|NOUN": 124.22, "art|NOUN": 123.8, "stödja|VERB": 123.76, "ond|ADJ": 123.18, "plan|NOUN": 52.0, "resa|NOUN": 122.43, "utom|ADP": 122.27, "hund|NOUN": 122.24, "syn|NOUN": 122.2, "glömma|VERB": 122.09, "avtal|NOUN": 121.92, "lek|NOUN": 121.7, "kul|ADJ": 121.6, "natt|NOUN": 121.51, "förändra|VERB": 121.43, "ange|VERB": 121.39, "någonting|PRON": 121.12, "förstås|ADV": 121.03, "individ|NOUN": 120.93, "älska|VERB": 120.93, "motion|NOUN": 120.87, "glad|ADJ": 120.57, "ned|PART": 120.5, "dator|NOUN": 120.28, "miljö|NOUN": 120.16, "ek|NOUN": 119.87, "åtminstone|ADV": 119.86, "presentera|VERB": 119.78, "stanna|VERB": 119.33, "byta|VERB": 119.29, "alternativ|NOUN": 118.94, "minut|NOUN": 118.87, "ingenting|PRON": 118.79, "uppleva|VERB": 118.65, "samla|VERB": 118.53, "svart|ADJ": 118.26, "bakgrund|NOUN": 118.12, "skott|NOUN": 118.07, "ö|NOUN": 118.02, "kärlek|NOUN": 118.0, "metod|NOUN": 117.61, "äldre|ADJ": 117.18, "säker|ADJ": 117.08, "borgare|NOUN": 117.01, "gud|NOUN": 116.98, "insats|NOUN": 116.63, "tysk|ADJ": 116.47, "kontroll|NOUN": 116.35, "lösa|VERB": 116.34, "kolla|VERB": 116.13, "fylla|VERB": 116.0, "bestämmelse|NOUN": 115.66, "ris|NOUN": 115.66, "drabba|VERB": 115.55, "nät|NOUN": 115.48, "teknik|NOUN": 115.08, "resurs|NOUN": 115.04, "försök|NOUN": 114.85, "fara|VERB": 114.82, "tjäna|VERB": 114.8, "argument|NOUN": 114.69, "behandla|VERB": 114.58, "ren|ADJ": 114.14, "fru|NOUN": 114.0, "sjuk|ADJ": 113.46, "istället för (el. i stället för)|ADP": 113.32, "våld|NOUN": 113.28, "utföra|VERB": 113.17, "ställning|NOUN": 113.06, "främst|ADV": 112.96, "räcka|VERB": 112.94, "bättre|ADV": 112.92, "fundera|VERB": 112.8, "visst|ADV": 112.62, "sommar|NOUN": 112.48, "rörelse|NOUN": 112.44, "kund|NOUN": 112.31, "villkor|NOUN": 112.19, "tillbaka (vardagl. tillbaks)|ADV": 112.16, "högt|ADV": 112.04, "president|NOUN": 111.99, "emellertid|ADV": 111.59, "händelse|NOUN": 111.44, "uppstå|VERB": 111.37, "acceptera|VERB": 111.33, "huvud|NOUN": 111.17, "sök|NOUN": 110.86, "snabb|ADJ": 110.8, "så kallad (förk. s.k., s k)|ADV": 110.51, "framför|ADP": 110.51, "ande|NOUN": 110.42, "bilda|VERB": 110.42, "orsak|NOUN": 110.42, "försvinna|VERB": 110.33, "fel|NOUN": 110.16, "innehåll|NOUN": 110.12, "natur|NOUN": 110.01, "begrepp|NOUN": 109.99, "för att|SCONJ": 109.47, "konflikt|NOUN": 109.19, "tack|INTJ": 108.87, "djur|NOUN": 108.73, "chans|NOUN": 108.16, "samtidigt som|SCONJ": 108.12, "demokratisk|ADJ": 107.94, "fel|ADV": 107.8, "läge|NOUN": 107.77, "sprida|VERB": 107.63, "växt|NOUN": 107.37, "förutom|ADP": 106.41, "i samband med|ADP": 106.3, "styck|NOUN": 106.25, "utskott|NOUN": 106.04, "muslim|NOUN": 105.98, "ordning|NOUN": 105.89, "uppdrag|NOUN": 105.87, "mark|NOUN": 105.63, "säkerhet|NOUN": 105.63, "linje|NOUN": 105.51, "bank|NOUN": 105.47, "önska|VERB": 105.47, "givetvis|ADV": 105.17, "studie|NOUN": 105.12, "fredag|NOUN": 104.7, "lärare|NOUN": 104.69, "statlig|ADJ": 104.45, "söndag|NOUN": 104.44, "fel|ADJ": 104.42, "speciellt|ADV": 104.35, "röd|ADJ": 104.34, "television (el. teve, tv)|NOUN": 104.3, "hot|NOUN": 104.27, "verk|NOUN": 104.0, "publicera|VERB": 103.98, "stund|NOUN": 103.98, "tillhöra|VERB": 103.16, "omfatta|VERB": 103.14, "material|NOUN": 102.94, "pelare|NOUN": 102.91, "hjärta|NOUN": 102.88, "knappast|ADV": 102.76, "befinna|VERB": 102.66, "part|NOUN": 102.65, "trevlig|ADJ": 102.64, "höst|NOUN": 102.61, "skilja|VERB": 102.57, "ens|ADV": 102.09, "förmåga|NOUN": 102.02, "döda|VERB": 101.92, "stånd|NOUN": 101.76, "peka|VERB": 101.73, "bedömning|NOUN": 101.49, "ringa|VERB": 101.34, "betrakta|VERB": 101.05, "by|NOUN": 100.93, "utifrån|ADP": 100.69, "brist|NOUN": 100.59, "hänga|VERB": 100.43, "tillräckligt|ADV": 100.4, "måndag|NOUN": 100.12, "aktuell|ADJ": 99.75, "någonsin (vardagl. nånsin)|ADV": 99.71, "tillåta|VERB": 99.66, "universitet|NOUN": 99.16, "konsekvens|NOUN": 99.15, "ställe|NOUN": 98.93, "hård|ADJ": 98.66, "majoritet|NOUN": 98.59, "domstol|NOUN": 98.49, "ordförande|NOUN": 98.46, "lördag|NOUN": 98.43, "låt|NOUN": 98.35, "herr|NOUN": 98.28, "sekvens|NOUN": 98.23, "förekomma|VERB": 98.18, "stoppa|VERB": 98.15, "nyhet|NOUN": 97.8, "journalist|NOUN": 97.73, "kris|NOUN": 97.59, "rycka|VERB": 97.44, "trycka|VERB": 97.44, "betydligt|ADV": 97.4, "kosta|VERB": 97.1, "band|NOUN": 97.09, "numera (el. numer)|ADV": 97.08, "tillstånd|NOUN": 97.07, "värd|ADJ": 97.06, "igen|PART": 96.98, "imorgon (el. i morgon)|ADV": 96.53, "klass|NOUN": 96.49, "uttrycka|VERB": 96.1, "slutsats|NOUN": 95.99, "global|ADJ": 95.78, "mitt|ADV": 95.61, "stol|NOUN": 95.52, "ytterligare|ADJ": 95.35, "effektiv|ADJ": 95.24, "resa|VERB": 95.16, "förbättra|VERB": 95.1, "rädda|VERB": 95.09, "list|NOUN": 94.89, "relation|NOUN": 94.81, "agera|VERB": 94.6, "central|ADJ": 94.56, "flera|PRON": 94.49, "undersökning|NOUN": 94.27, "uppnå|VERB": 94.18, "krona (förk. kr.)|NOUN": 94.15, "perspektiv|NOUN": 94.04, "plötsligt|ADV": 93.95, "naturlig|ADJ": 93.87, "ålder|NOUN": 93.87, "process|NOUN": 93.76, "uttryck|NOUN": 93.7, "lista|NOUN": 93.66, "allra|ADV": 93.57, "sökning|NOUN": 93.56, "ökning|NOUN": 93.56, "därför att|SCONJ": 93.55, "rysk|ADJ": 93.55, "jämföra (förk. jfr)|VERB": 93.52, "tills|SCONJ": 93.48, "intresserad|ADJ": 93.21, "totalt|ADV": 92.97, "hantera|VERB": 92.87, "förvänta|VERB": 92.79, "medel|NOUN": 92.73, "vika|VERB": 92.39, "döma|VERB": 92.38, "besöka|VERB": 92.36, "hem|NOUN": 92.26, "var|ADV": 92.16, "täcka|VERB": 92.1, "borgerlig|ADJ": 92.09, "inleda|VERB": 92.09, "helg|NOUN": 92.06, "undvika|VERB": 92.02, "ryck|NOUN": 91.76, "tryck|NOUN": 91.76, "tydligen|ADV": 91.69, "aktiv|ADJ": 91.62, "höja|VERB": 91.58, "pappa|NOUN": 91.48, "varkeneller|CCONJ": 91.32, "religiös|ADJ": 91.15, "råka|VERB": 91.0, "verklig|ADJ": 90.87, "rent|ADV": 90.85, "fantastisk|ADJ": 90.78, "grundläggande|ADJ": 90.73, "upptäcka|VERB": 90.72, "erkänna|VERB": 90.67, "helig|ADJ": 90.59, "lön|NOUN": 90.42, "historisk|ADJ": 90.34, "rest|NOUN": 90.27, "halv|ADJ": 90.13, "andel|NOUN": 90.06, "besök|NOUN": 90.06, "teknisk|ADJ": 90.04, "kasta|VERB": 89.78, "hemsida|NOUN": 89.75, "bedöma|VERB": 89.72, "torsdag|NOUN": 89.68, "tillväxt|NOUN": 89.64, "läsare|NOUN": 89.59, "forskare|NOUN": 89.52, "bidrag|NOUN": 89.28, "onsdag|NOUN": 89.16, "vilja|NOUN": 89.16, "sol|NOUN": 89.1, "inte minst|ADV": 89.08, "analys|NOUN": 88.93, "ovan|ADV": 88.85, "lagstiftning|NOUN": 88.83, "militär|ADJ": 88.82, "toppa|VERB": 88.72, "sort|NOUN": 88.57, "fördel|NOUN": 88.33, "skydda|VERB": 88.3, "nyttja|VERB": 88.29, "utnyttja|VERB": 88.29, "teori|NOUN": 88.16, "fransk|ADJ": 88.02, "pågå|VERB": 87.99, "samling|NOUN": 87.94, "flertal|NOUN": 87.89, "snarare|ADV": 87.88, "försvara|VERB": 87.72, "modell|NOUN": 87.56, "skön|ADJ": 87.52, "vapen|NOUN": 87.52, "således|ADV": 87.49, "förening|NOUN": 87.48, "lyfta|VERB": 87.39, "eftermiddag (förk. em.)|NOUN": 87.36, "soldat|NOUN": 87.29, "märka|VERB": 87.24, "gemenskap|NOUN": 87.17, "ösa|VERB": 87.12, "fast|CCONJ": 87.09, "styrka|NOUN": 86.87, "ersätta|VERB": 86.51, "kille|NOUN": 86.47, "vård|NOUN": 86.44, "fullt|ADV": 86.4, "ägna|VERB": 86.39, "oavsett|ADP": 86.16, "poäng|NOUN": 86.13, "satsa|VERB": 86.11, "moderat|NOUN": 86.02, "rida|VERB": 85.96, "jo|INTJ": 85.95, "tisdag|NOUN": 85.94, "död|ADJ": 85.9, "allmänt|ADV": 85.48, "avsluta|VERB": 85.39, "sova|VERB": 85.26, "inne|ADV": 85.1, "flicka|NOUN": 85.02, "sedan (vardagl. sen)|SCONJ": 84.79, "total|ADJ": 84.78, "allvarlig|ADJ": 84.74, "fram|ADV": 84.73, "ljus|NOUN": 84.31, "sjukdom|NOUN": 84.27, "unge|NOUN": 84.16, "i form av|ADP": 84.01, "vikt|NOUN": 83.95, "rik|ADJ": 83.8, "region|NOUN": 83.76, "samtal|NOUN": 83.69, "negativ|ADJ": 83.54, "mycket|PRON": 83.53, "i år|ADV": 83.52, "igång|PART": 83.49, "vändning|NOUN": 83.42, "antingeneller|CCONJ": 83.19, "föda|VERB": 83.1, "åter|ADV": 83.06, "arbetare|NOUN": 83.02, "skjuta|VERB": 83.01, "tradition|NOUN": 82.91, "hämta|VERB": 82.84, "församling|NOUN": 82.73, "hav|NOUN": 82.66, "energi|NOUN": 82.37, "bred|ADJ": 82.28, "vad gäller|ADP": 82.23, "fast|PART": 82.22, "påpeka|VERB": 82.21, "bättra|VERB": 82.19, "skaffa|VERB": 82.09, "utgå|VERB": 82.08, "samtlig|ADJ": 81.95, "stärka|VERB": 81.95, "läkare|NOUN": 81.81, "fattig|ADJ": 81.56, "grepp|NOUN": 81.5, "hej|INTJ": 81.45, "utsätta|VERB": 81.45, "spännande|ADJ": 81.2, "fort|ADV": 81.07, "sikt|NOUN": 81.06, "revolution|NOUN": 81.03, "brev|NOUN": 80.95, "personal|NOUN": 80.84, "skada|NOUN": 80.74, "illa|ADV": 80.73, "kämpa|VERB": 80.69, "alltför|ADV": 80.65, "tecken|NOUN": 80.61, "siffra|NOUN": 80.59, "tydligt|ADV": 80.52, "än (el. ännu)|ADV": 80.5, "hårt|ADV": 80.46, "absolut|ADV": 80.27, "eka|VERB": 80.26, "engelsk|ADJ": 80.2, "praktik|NOUN": 79.79, "förmodligen|ADV": 79.75, "hoppa|VERB": 79.72, "morgon|NOUN": 79.54, "tjej|NOUN": 79.44, "konstig|ADJ": 79.43, "union|NOUN": 79.39, "kommande|ADJ": 79.27, "avgöra|VERB": 79.23, "chef|NOUN": 79.17, "vis|NOUN": 79.11, "strid|NOUN": 78.98, "sända|VERB": 78.93, "missa|VERB": 78.88, "bedriva|VERB": 78.64, "etcetera (el. et cetera, förk. etc.)|ADV": 78.45, "anföra|VERB": 78.34, "varm|ADJ": 78.22, "hit|ADV": 78.19, "berättelse|NOUN": 78.05, "produktion|NOUN": 77.86, "kapitel (förk. kap.)|NOUN": 77.76, "hindra|VERB": 77.58, "konst|NOUN": 77.53, "speciell|ADJ": 77.45, "allvar|NOUN": 77.42, "grön|ADJ": 77.31, "vår|NOUN": 77.26, "meddela|VERB": 77.16, "omöjlig|ADJ": 77.05, "tillämpa|VERB": 77.02, "skydd|NOUN": 76.99, "hittills|ADV": 76.96, "sällan|ADV": 76.95, "position|NOUN": 76.89, "behandling|NOUN": 76.64, "omfattande|ADJ": 76.54, "skog|NOUN": 76.52, "kritisera|VERB": 76.46, "förklaring|NOUN": 76.39, "springa|VERB": 76.39, "oerhört|ADV": 76.26, "uppfatta|VERB": 76.24, "foto|NOUN": 76.14, "islam|NOUN": 76.13, "stänga|VERB": 76.1, "aning|NOUN": 76.09, "försvar|NOUN": 76.08, "meter|NOUN": 76.04, "evolution|NOUN": 75.98, "funktion|NOUN": 75.88, "dotter|NOUN": 75.82, "värdering|NOUN": 75.62, "råda|VERB": 75.56, "ersättning|NOUN": 75.51, "slippa|VERB": 75.51, "självklart|ADV": 75.31, "lämplig|ADJ": 75.27, "ting|NOUN": 75.13, "minne|NOUN": 75.11, "strategi|NOUN": 75.1, "dyka|VERB": 75.09, "orka|VERB": 75.09, "kontrollera|VERB": 74.97, "planera|VERB": 74.86, "färg|NOUN": 74.81, "lova|VERB": 74.62, "citera|VERB": 74.41, "finansiell|ADJ": 74.34, "ständigt|ADV": 74.22, "spår|NOUN": 74.17, "kall|ADJ": 74.14, "vuxen|ADJ": 74.07, "allians|NOUN": 74.06, "faktor|NOUN": 73.95, "kvalitet (el. kvalité)|NOUN": 73.93, "upp|ADV": 73.89, "utländsk|ADJ": 73.89, "svag|ADJ": 73.87, "sköta|VERB": 73.72, "vägra|VERB": 73.64, "rike|NOUN": 73.5, "framgå|VERB": 73.41, "judisk|ADJ": 73.26, "studera|VERB": 73.17, "farlig|ADJ": 73.07, "framgång|NOUN": 73.07, "tolka|VERB": 73.02, "billig|ADJ": 73.02, "iväg|PART": 72.74, "student|NOUN": 72.69, "och så vidare (förk. o.s.v., osv.)|ADV": 72.62, "visserligen|ADV": 72.58, "vara|NOUN": 72.57, "undantag|NOUN": 72.4, "tillgänglig|ADJ": 72.31, "enorm|ADJ": 72.24, "behålla|VERB": 72.2, "dricka|VERB": 72.16, "aktion|NOUN": 72.14, "bry sig|VERB": 72.13, "relativt|ADV": 72.06, "tung|ADJ": 72.04, "arbetsgivare|NOUN": 71.89, "med hjälp av|ADP": 71.84, "tvärtom (el. tvärt om)|ADV": 71.67, "notera|VERB": 71.48, "nation|NOUN": 71.44, "sänka|VERB": 71.42, "ärende|NOUN": 71.39, "givare|NOUN": 71.09, "kull|NOUN": 71.03, "nyligen|ADV": 71.03, "rättelse|NOUN": 71.0, "delvis|ADV": 70.94, "medföra|VERB": 70.92, "ifrågasätta|VERB": 70.79, "för övrigt|ADV": 70.76, "län|NOUN": 70.61, "gata|NOUN": 70.48, "medveten|ADJ": 70.44, "serie|NOUN": 70.44, "rimlig|ADJ": 70.42, "ty|CCONJ": 70.38, "invandrare|NOUN": 70.38, "dörr|NOUN": 70.02, "direktiv|NOUN": 69.99, "stiga|VERB": 69.91, "tiga|VERB": 69.91, "fot|NOUN": 69.9, "begränsad|ADJ": 69.9, "vag|ADJ": 69.88, "äntligen|ADV": 69.88, "vänster|ADJ": 69.77, "ner (el. ned)|ADV": 69.65, "väcka|VERB": 69.65, "leta|VERB": 69.52, "häst|NOUN": 69.47, "kategori|NOUN": 69.47, "brittisk|ADJ": 69.43, "följd|NOUN": 69.24, "ed|NOUN": 69.22, "fred|NOUN": 69.22, "traditionell|ADJ": 69.22, "användning|NOUN": 69.21, "riskera|VERB": 69.16, "tappa|VERB": 69.16, "inkomst|NOUN": 69.04, "nöjd|ADJ": 69.02, "kläder|NOUN": 69.0, "spara|VERB": 68.81, "styrelse|NOUN": 68.79, "intervju|NOUN": 68.72, "starkt|ADV": 68.69, "slutligen|ADV": 68.46, "bit|NOUN": 68.3, "muslimsk|ADJ": 68.24, "vetenskaplig|ADJ": 68.23, "överens|ADV": 67.86, "framtida|ADJ": 67.84, "bevis|NOUN": 67.69, "fast|ADJ": 67.58, "sexuell|ADJ": 67.49, "exakt|ADV": 67.27, "arbetsmarknad|NOUN": 67.26, "underbar|ADJ": 67.23, "post|NOUN": 67.02, "extra|ADJ": 66.9, "offer|NOUN": 66.85, "sektor|NOUN": 66.75, "vinst|NOUN": 66.65, "England|PROPN": 66.6, "inflytande|NOUN": 66.6, "budskap|NOUN": 66.59, "klicka|VERB": 66.58, "tips|NOUN": 66.37, "världskrig|NOUN": 66.36, "med tanke på|ADP": 66.31, "självklar|ADJ": 66.24, "båt|NOUN": 66.17, "borta|ADV": 66.14, "regional|ADJ": 66.06, "framåt|ADV": 66.04, "karaktär|NOUN": 66.0, "skiva|NOUN": 66.0, "omkring|ADV": 65.97, "ansikte|NOUN": 65.96, "i början|ADP": 65.88, "aktivitet|NOUN": 65.76, "ost|NOUN": 65.67, "fängelse|NOUN": 65.6, "motsvarande|ADJ": 65.56, "synas|VERB": 65.54, "mor (el. moder, vardagl. morsa) |NOUN": 65.46, "an|PART": 65.44, "samman|PART": 65.44, "ända|ADV": 65.38, "ledamot|NOUN": 65.34, "i enlighet med|ADP": 65.2, "civil|ADJ": 65.17, "uppenbar|ADJ": 65.12, "skull|NOUN": 65.07, "arbetslöshet|NOUN": 65.0, "fysisk|ADJ": 64.96, "generation|NOUN": 64.92, "återigen|ADV": 64.84, "djup|ADJ": 64.61, "initiativ|NOUN": 64.56, "fastställa|VERB": 64.47, "parlament|NOUN": 64.38, "säsong|NOUN": 64.38, "levande|ADJ": 64.27, "tacka|VERB": 64.24, "hota|VERB": 64.07, "tusentals|ADV": 64.02, "eventuell|ADJ": 64.0, "pojke|NOUN": 63.91, "version|NOUN": 63.9, "existera|VERB": 63.72, "trött|ADJ": 63.63, "himmel|NOUN": 63.39, "reaktion|NOUN": 63.39, "dyr|ADJ": 63.35, "normal|ADJ": 63.27, "rikta|VERB": 63.25, "kurs|NOUN": 63.24, "påstående|NOUN": 63.24, "märklig|ADJ": 63.17, "öst|NOUN": 63.12, "affär|NOUN": 63.08, "tidigt|ADV": 62.99, "upplevelse|NOUN": 62.97, "riktning|NOUN": 62.93, "vetenskap|NOUN": 62.83, "avsnitt|NOUN": 62.81, "handel|NOUN": 62.81, "sträckning|NOUN": 62.79, "locka|VERB": 62.67, "redovisa|VERB": 62.59, "uttalande|NOUN": 62.58, "respektive|CCONJ": 62.53, "para|VERB": 62.49, "störa|VERB": 62.42, "ihåg|PART": 62.4, "någonstans (vardagl. nånstans)|ADV": 62.31, "respekt|NOUN": 62.24, "rapportera|VERB": 62.23, "knappt|ADV": 62.21, "direkt|ADJ": 62.17, "enkelt|ADV": 62.17, "omständighet|NOUN": 62.09, "hänsyn|NOUN": 62.05, "ikväll (el. i kväll)|ADV": 62.03, "begära|VERB": 61.92, "rubrik|NOUN": 61.88, "producera|VERB": 61.86, "utsträckning|NOUN": 61.82, "anonym|ADJ": 61.81, "begå|VERB": 61.74, "bar|ADJ": 61.59, "institution|NOUN": 61.59, "förstöra|VERB": 61.58, "boll|NOUN": 61.53, "grunda|VERB": 61.49, "förbi|ADP": 61.34, "luft|NOUN": 61.33, "industri|NOUN": 61.23, "tåg|NOUN": 61.07, "skada|VERB": 61.02, "nordisk|ADJ": 60.93, "uppfylla|VERB": 60.84, "akta|VERB": 60.82, "förhandling|NOUN": 60.69, "syfta|VERB": 60.6, "bror (el. broder, vardagl. brorsa)|NOUN": 60.45, "byggnad|NOUN": 60.45, "hälft|NOUN": 60.43, "skrift|NOUN": 60.43, "ansvarig|ADJ": 60.34, "allmänhet|NOUN": 60.26, "orsaka|VERB": 60.24, "i slutet|ADP": 60.23, "israelisk|ADJ": 60.2, "drygt|ADV": 60.1, "lever|NOUN": 60.09, "bloggare|NOUN": 60.07, "tävling|NOUN": 59.87, "kommunikation|NOUN": 59.79, "kritisk|ADJ": 59.66, "plocka|VERB": 59.59, "patient|NOUN": 59.58, "sjunga|VERB": 59.53, "vakna|VERB": 59.51, "hälsa|NOUN": 59.45, "piratparti|NOUN": 59.45, "centrum|NOUN": 59.43, "otroligt|ADV": 59.42, "roligt|ADV": 59.42, "mörk|ADJ": 59.31, "träna|VERB": 59.09, "bord|NOUN": 59.07, "förrän|SCONJ": 59.06, "dansk|ADJ": 59.05, "vidta|VERB": 59.02, "reda|NOUN": 59.02, "mana|VERB": 58.88, "väljare|NOUN": 58.84, "uppmana|VERB": 58.76, "publik|NOUN": 58.71, "lida|VERB": 58.6, "motstånd|NOUN": 58.6, "lägenhet|NOUN": 58.56, "vänsterparti|NOUN": 58.46, "rädd|ADJ": 58.45, "användare|NOUN": 58.35, "inre|ADJ": 58.31, "avslöja|VERB": 58.29, "fiende|NOUN": 58.26, "lopp|NOUN": 58.2, "återvända|VERB": 58.17, "utmaning|NOUN": 58.16, "hopp|NOUN": 58.14, "konkurrens|NOUN": 58.14, "dröm|NOUN": 58.07, "detalj|NOUN": 58.03, "nedan|ADV": 57.98, "placera|VERB": 57.94, "litteratur|NOUN": 57.85, "ana|VERB": 57.79, "inställning|NOUN": 57.78, "armé|NOUN": 57.72, "lös|ADJ": 57.71, "pröva|VERB": 57.64, "egenskap|NOUN": 57.61, "rekommendera|VERB": 57.61, "liberal|ADJ": 57.58, "synpunkt|NOUN": 57.51, "undan|ADP": 57.5, "angående|ADP": 57.49, "unik|ADJ": 57.46, "präst|NOUN": 57.44, "webbplats|NOUN": 57.41, "bostad|NOUN": 57.37, "vardag|NOUN": 57.37, "gratis|ADV": 57.31, "återkomma|VERB": 57.2, "bevisa|VERB": 57.17, "anställd|NOUN": 57.15, "förbjuda|VERB": 57.13, "uttala|VERB": 57.08, "investering|NOUN": 57.01, "fira|VERB": 56.93, "försäljning|NOUN": 56.93, "populär|ADJ": 56.93, "klubb|NOUN": 56.9, "citat|NOUN": 56.87, "palestinier|NOUN": 56.84, "utrymme|NOUN": 56.83, "förr|ADV": 56.75, "svårt|ADV": 56.72, "stark|ADJ": 56.58, "påminna|VERB": 56.57, "aktör|NOUN": 56.53, "klassisk|ADJ": 56.38, "omkring|ADP": 56.37, "fokus|NOUN": 56.32, "officiell|ADJ": 56.31, "beröra|VERB": 56.26, "palestinsk|ADJ": 56.26, "ägare|NOUN": 56.2, "kapital|NOUN": 56.03, "relevant|ADJ": 56.02, "minister|NOUN": 55.85, "anpassa|VERB": 55.79, "glädje|NOUN": 55.79, "titel|NOUN": 55.79, "något|ADV": 55.74, "utgångspunkt|NOUN": 55.74, "nätverk|NOUN": 55.73, "scen|NOUN": 55.67, "nytta|NOUN": 55.62, "hållbar|ADJ": 55.61, "begränsa|VERB": 55.6, "sikte|NOUN": 55.52, "snygg|ADJ": 55.44, "kvinnlig|ADJ": 55.42, "som vanligt|ADV": 55.42, "avstånd|NOUN": 55.37, "fly|VERB": 55.32, "betydande|ADJ": 55.32, "skyldig|ADJ": 55.31, "i övrigt|ADV": 55.3, "inflation|NOUN": 55.13, "ben|NOUN": 55.11, "definition|NOUN": 54.94, "uppmärksamhet|NOUN": 54.9, "ladda|VERB": 54.89, "jul|NOUN": 54.78, "dåligt|ADV": 54.56, "kommunal|ADJ": 54.45, "passera|VERB": 54.39, "herre|NOUN": 54.34, "i fråga om|ADP": 54.28, "klimat|NOUN": 54.24, "var|PRON": 54.15, "topp|NOUN": 54.11, "troligen|ADV": 54.11, "kompis|NOUN": 53.95, "främja|VERB": 53.95, "landsting|NOUN": 53.95, "undersöka|VERB": 53.89, "kilometer (förk. km)|NOUN": 53.72, "reform|NOUN": 53.71, "testa|VERB": 53.66, "konkret|ADJ": 53.61, "rakt|ADV": 53.53, "uppenbarligen|ADV": 53.53, "desto|ADV": 53.5, "socialdemokratisk|ADJ": 53.5, "trupp|NOUN": 53.44, "vart|ADV": 53.43, "seger|NOUN": 53.38, "centerparti|NOUN": 53.37, "förlust|NOUN": 53.3, "själ|NOUN": 53.26, "öde|NOUN": 53.22, "mord|NOUN": 53.2, "dokument|NOUN": 53.17, "upphöra|VERB": 53.15, "folkparti|NOUN": 53.14, "kraftigt|ADV": 53.14, "middag|NOUN": 53.1, "reagera|VERB": 53.1, "hjärna|NOUN": 53.02, "kulturell|ADJ": 53.02, "södra|ADJ": 53.02, "fast|SCONJ": 53.01, "förtroende|NOUN": 52.99, "förordning|NOUN": 52.95, "upphovsrätt|NOUN": 52.95, "skuld|NOUN": 52.87, "professor|NOUN": 52.61, "inklusive|ADP": 52.53, "beskrivning|NOUN": 52.51, "lycka|NOUN": 52.51, "skrivning|NOUN": 52.51, "yrkande|NOUN": 52.51, "kär|ADJ": 52.5, "äng|NOUN": 52.49, "hänvisa|VERB": 52.38, "buss|NOUN": 52.35, "norra|ADJ": 52.24, "fullständigt|ADV": 52.21, "make|NOUN": 52.21, "antagligen|ADV": 52.05, "stil|NOUN": 51.78, "förbund|NOUN": 51.74, "tolkning|NOUN": 51.7, "utöver|ADP": 51.6, "syster (vardagl. syrra)|NOUN": 51.59, "berg|NOUN": 51.57, "motståndare|NOUN": 51.53, "höger|ADJ": 51.47, "praktisk|ADJ": 51.45, "beteende|NOUN": 51.29, "bud|NOUN": 51.28, "träning|NOUN": 51.25, "vare sig|CCONJ": 51.25, "äktenskap|NOUN": 51.11, "grov|ADJ": 51.04, "uppe|ADV": 50.95, "inslag|NOUN": 50.92, "förhindra|VERB": 50.9, "delning|NOUN": 50.82, "kapitalism|NOUN": 50.81, "bilaga|NOUN": 50.76, "tom|ADJ": 50.74, "invånare|NOUN": 50.64, "struktur|NOUN": 50.56, "politiskt|ADV": 50.53, "sjukhus|NOUN": 50.51, "mer eller mindre|ADV": 50.5, "främsta|ADJ": 50.47, "djupt|ADV": 50.43, "visning|NOUN": 50.3, "korrekt|ADJ": 50.24, "bäst|ADV": 50.24, "gentemot|ADP": 50.23, "tack vare|ADP": 50.23, "aspekt|NOUN": 50.22, "godkänna|VERB": 50.2, "felaktig|ADJ": 50.17, "dialog|NOUN": 50.17, "oro|NOUN": 50.14, "vägg|NOUN": 50.14, "kinesisk|ADJ": 50.13, "ständig|ADJ": 50.11, "tema|NOUN": 50.11, "helhet|NOUN": 50.05, "satsning|NOUN": 50.02, "statistik|NOUN": 50.0, "beräkna|VERB": 49.99, "resonemang|NOUN": 49.97, "förbud|NOUN": 49.95, "dollar|NOUN": 49.94, "längs|ADP": 49.8, "fixa|VERB": 49.79, "kollega|NOUN": 49.68, "inträffa|VERB": 49.66, "sjukvård|NOUN": 49.6, "överleva|VERB": 49.51, "sannolikt|ADV": 49.49, "i första hand|ADV": 49.48, "meddelande|NOUN": 49.48, "näringsliv|NOUN": 49.43, "låna|VERB": 49.26, "förståelse|NOUN": 49.23, "möjligen|ADV": 49.17, "fisk|NOUN": 49.17, "konsument|NOUN": 49.13, "framhålla|VERB": 49.07, "storlek|NOUN": 49.07, "telefon|NOUN": 48.95, "kön|NOUN": 48.94, "slut|PART": 48.93, "laga|VERB": 48.7, "roman|NOUN": 48.7, "lån|NOUN": 48.68, "likna|VERB": 48.67, "lita|VERB": 48.62, "säng|NOUN": 48.59, "rädsla|NOUN": 48.56, "övertygad|ADJ": 48.55, "skit|NOUN": 48.52, "tänkande|NOUN": 48.51, "arm|NOUN": 48.45, "bruk|NOUN": 48.4, "radio|NOUN": 48.33, "granska|VERB": 48.31, "i synnerhet|ADV": 48.31, "bekräfta|VERB": 48.27, "väder|NOUN": 48.25, "hinder|NOUN": 48.24, "förut|ADV": 48.23, "personligen|ADV": 48.21, "bana|NOUN": 48.15, "reklam|NOUN": 48.04, "trafik|NOUN": 48.01, "ärlig|ADJ": 47.97, "allting|PRON": 47.95, "artist|NOUN": 47.95, "bröd|NOUN": 47.92, "huruvida|SCONJ": 47.92, "utsatt|ADJ": 47.92, "butik|NOUN": 47.83, "ytterst|ADV": 47.74, "förbli|VERB": 47.73, "tråkig|ADJ": 47.67, "hemlig|ADJ": 47.62, "andlig|ADJ": 47.6, "beträffande|ADP": 47.59, "vänster|NOUN": 47.58, "fartyg|NOUN": 47.47, "flyga|VERB": 47.45, "gifta|VERB": 47.43, "snäll|ADJ": 47.36, "ränta|NOUN": 47.34, "proposition|NOUN": 47.31, "svårighet|NOUN": 47.24, "fart|NOUN": 47.21, "tant|NOUN": 47.2, "berörd|ADJ": 47.13, "avsikt|NOUN": 47.12, "frisk|ADJ": 47.12, "opposition|NOUN": 47.11, "härlig|ADJ": 47.1, "intryck|NOUN": 47.0, "visa|NOUN": 46.94, "duktig|ADJ": 46.87, "ideologi|NOUN": 46.83, "representant|NOUN": 46.77, "tack|NOUN": 46.74, "engagemang|NOUN": 46.69, "finsk|ADJ": 46.66, "bekant|ADJ": 46.6, "överallt|ADV": 46.57, "gäng|NOUN": 46.56, "träda|VERB": 46.56, "sjunka|VERB": 46.55, "föremål|NOUN": 46.54, "vad|ADV": 46.51, "attack|NOUN": 46.49, "falsk|ADJ": 46.49, "representera|VERB": 46.46, "miljöparti|NOUN": 46.41, "avgift|NOUN": 46.38, "normalt|ADV": 46.36, "motsvara|VERB": 46.25, "i allmänhet|ADV": 46.2, "översättning|NOUN": 46.2, "seriös|ADJ": 46.16, "omedelbart|ADV": 46.15, "kraftig|ADJ": 46.13, "uppskatta|VERB": 46.1, "kommitté|NOUN": 46.0, "blanda|VERB": 45.98, "blod|NOUN": 45.98, "högskola|NOUN": 45.98, "fritt|ADV": 45.9, "integritet|NOUN": 45.9, "hår|NOUN": 45.86, "organ|NOUN": 45.79, "lycklig|ADJ": 45.77, "misstag|NOUN": 45.74, "kvar|ADV": 45.69, "träd|NOUN": 45.68, "tak|NOUN": 45.67, "straff|NOUN": 45.66, "perfekt|ADJ": 45.65, "överenskommelse|NOUN": 45.61, "kampanj|NOUN": 45.59, "grej|NOUN": 45.58, "åstadkomma|VERB": 45.57, "budget|NOUN": 45.56, "rygg|NOUN": 45.55, "gott|ADV": 45.5, "press|NOUN": 45.45, "digital|ADJ": 45.42, "framstå|VERB": 45.4, "verktyg|NOUN": 45.4, "beroende på|ADP": 45.39, "betyg|NOUN": 45.28, "detsamma|PRON": 45.26, "start|NOUN": 45.17, "leverera|VERB": 45.14, "kompetens|NOUN": 45.13, "var och en|PRON": 45.08, "långsiktig|ADJ": 44.96, "vinter|NOUN": 44.95, "gripa|VERB": 44.94, "skyldighet|NOUN": 44.81, "evig|ADJ": 44.78, "företrädare|NOUN": 44.73, "etnisk|ADJ": 44.59, "med andra ord|ADV": 44.51, "njuta|VERB": 44.46, "posta|VERB": 44.39, "runda|VERB": 44.38, "för|CCONJ": 44.36, "bereda|VERB": 44.28, "uppmärksamma|VERB": 44.27, "arbetslös|ADJ": 44.2, "yta|NOUN": 44.18, "skratta|VERB": 44.04, "underlätta|VERB": 44.04, "föreligga|VERB": 43.98, "tillämpning|NOUN": 43.98, "garantera|VERB": 43.97, "jakt|NOUN": 43.94, "utse|VERB": 43.93, "blick|NOUN": 43.86, "svenska|NOUN": 43.74, "konferens|NOUN": 43.68, "framföra|VERB": 43.66, "runt|ADV": 43.65, "specifik|ADJ": 43.64, "varg|NOUN": 43.6, "kanal|NOUN": 43.59, "klok|ADJ": 43.53, "regim|NOUN": 43.51, "utöva|VERB": 43.51, "fokusera|VERB": 43.48, "belopp|NOUN": 43.46, "bransch|NOUN": 43.46, "sekund|NOUN": 43.43, "reda|VERB": 43.42, "torde|AUX": 43.35, "färdig|ADJ": 43.33, "ordna|VERB": 43.33, "närma|VERB": 43.31, "vind|NOUN": 43.29, "gård|NOUN": 43.28, "mitt|NOUN": 43.27, "framgångsrik|ADJ": 43.21, "identitet|NOUN": 43.18, "sång|NOUN": 43.18, "närma sig|VERB": 43.14, "skrika|VERB": 43.14, "tidpunkt|NOUN": 43.12, "avskaffa|VERB": 43.11, "samband|NOUN": 43.1, "lugn|ADJ": 43.08, "uppge|VERB": 43.08, "deltagare|NOUN": 43.07, "ursprung|NOUN": 43.07, "bestämd|ADJ": 43.06, "insikt|NOUN": 43.05, "forum|NOUN": 43.03, "kort|NOUN": 43.02, "statsminister|NOUN": 42.87, "annorlunda|ADJ": 42.85, "definiera|VERB": 42.8, "fönster|NOUN": 42.75, "get|NOUN": 42.71, "likhet|NOUN": 42.68, "ljud|NOUN": 42.67, "beställa|VERB": 42.48, "synd|NOUN": 42.46, "papper|NOUN": 42.43, "fara|NOUN": 42.39, "definitivt|ADV": 42.38, "omfattning|NOUN": 42.37, "bevara|VERB": 42.29, "väga|VERB": 42.23, "fenomen|NOUN": 42.2, "riktlinje|NOUN": 42.17, "profet|NOUN": 42.16, "decennium|NOUN": 42.15, "i stort sett|ADV": 42.1, "inriktning|NOUN": 42.05, "misslyckas|VERB": 42.04, "ram|NOUN": 42.04, "finansiera|VERB": 42.03, "hotell|NOUN": 42.0, "kristendom|NOUN": 42.0, "dess|ADV": 41.98, "i förhållande till|ADP": 41.87, "klaga|VERB": 41.87, "skatta|VERB": 41.87, "upprätta|VERB": 41.86, "förhoppningsvis|ADV": 41.58, "gynna|VERB": 41.53, "ifall|SCONJ": 41.43, "oberoende|ADJ": 41.42, "leka|VERB": 41.37, "märke|NOUN": 41.31, "snö|NOUN": 41.31, "upprepa|VERB": 41.31, "undervisning|NOUN": 41.29, "kött|NOUN": 41.19, "förutsätta|VERB": 41.16, "replik|NOUN": 41.12, "koppling|NOUN": 41.1, "snitt|NOUN": 41.04, "engelska|NOUN": 41.03, "överhuvudtaget|ADV": 41.0, "sysselsättning|NOUN": 40.97, "besked|NOUN": 40.96, "lätta|VERB": 40.92, "oavsett|ADV": 40.87, "avseende|NOUN": 40.83, "okänd|ADJ": 40.81, "katolsk|ADJ": 40.79, "ropa|VERB": 40.76, "bekämpa|VERB": 40.74, "synd|ADV": 40.74, "genast|ADV": 40.7, "sjö|NOUN": 40.7, "så småningom (el. småningom)|ADV": 40.7, "logisk|ADJ": 40.69, "inom ramen för|ADP": 40.67, "kaffe|NOUN": 40.67, "förstärka|VERB": 40.65, "euro|NOUN": 40.64, "mänsklighet|NOUN": 40.59, "nere|ADV": 40.57, "betona|VERB": 40.53, "expert|NOUN": 40.48, "fildelning|NOUN": 40.41, "olja|NOUN": 40.38, "förbereda|VERB": 40.33, "förfarande|NOUN": 40.3, "trygghet|NOUN": 40.26, "konstnär|NOUN": 40.2, "i själva verket|ADV": 40.15, "norsk|ADJ": 40.15, "i fråga (el. ifråga)|ADV": 40.14, "stjärna|NOUN": 40.12, "tyg|NOUN": 40.09, "läsning|NOUN": 40.01, "blå|ADJ": 40.0, "fotboll|NOUN": 40.0, "flykting|NOUN": 39.98, "koppla|VERB": 39.9, "forma|VERB": 39.88, "bibel|NOUN": 39.87, "förresten|ADV": 39.86, "samarbeta|VERB": 39.84, "slänga|VERB": 39.82, "ögonblick|NOUN": 39.81, "neka|VERB": 39.75, "extra|ADV": 39.67, "arbetsplats|NOUN": 39.66, "lokal|NOUN": 39.58, "summa|NOUN": 39.56, "tillräcklig|ADJ": 39.49, "äcklig|ADJ": 39.49, "tona|VERB": 39.44, "tendens|NOUN": 39.43, "på så sätt|ADV": 39.33, "restaurang|NOUN": 39.29, "återstå|VERB": 39.29, "vila|VERB": 39.26, "extremt|ADV": 39.25, "kamera|NOUN": 39.24, "självständig|ADJ": 39.17, "socialistisk|ADJ": 39.15, "framställa|VERB": 39.04, "ända (el. ände)|NOUN": 39.0, "mångfald|NOUN": 38.97, "strand|NOUN": 38.97, "pension|NOUN": 38.96, "hem|ADV": 38.95, "diskriminering|NOUN": 38.94, "misstänka|VERB": 38.94, "utsläpp|NOUN": 38.92, "logga|VERB": 38.85, "medicin|NOUN": 38.84, "sport|NOUN": 38.76, "rättvisa|NOUN": 38.74, "eld|NOUN": 38.73, "individuell|ADJ": 38.72, "därifrån|ADV": 38.64, "ifrån|ADV": 38.64, "yttre|ADJ": 38.53, "arabisk|ADJ": 38.42, "erhålla|VERB": 38.41, "moralisk|ADJ": 38.41, "revolutionär|ADJ": 38.4, "egendom|NOUN": 38.38, "köp|NOUN": 38.33, "välfärd|NOUN": 38.32, "sticka|VERB": 38.31, "mäta|VERB": 38.3, "helvete|NOUN": 38.27, "tuff|ADJ": 38.27, "jordbruk|NOUN": 38.26, "sällskap|NOUN": 38.25, "medverka|VERB": 38.2, "arbetstagare|NOUN": 38.17, "fånga|VERB": 38.16, "blogga|VERB": 38.15, "terrorism|NOUN": 38.13, "fest|NOUN": 38.12, "ordentligt|ADV": 38.12, "väst|NOUN": 38.1, "sajt|NOUN": 38.08, "prova|VERB": 38.07, "prägla|VERB": 38.03, "dum|ADJ": 38.02, "övning|NOUN": 37.99, "jobbig|ADJ": 37.96, "måla|VERB": 37.96, "vin|NOUN": 37.91, "identifiera|VERB": 37.89, "rasism|NOUN": 37.84, "ståndpunkt|NOUN": 37.84, "granne|NOUN": 37.82, "rang|NOUN": 37.81, "resultera|VERB": 37.79, "karriär|NOUN": 37.72, "trend|NOUN": 37.69, "kontor|NOUN": 37.63, "jaga|VERB": 37.6, "yttrandefrihet|NOUN": 37.57, "fortsättning|NOUN": 37.46, "diverse|ADJ": 37.46, "stöta|VERB": 37.45, "förneka|VERB": 37.44, "väsentlig|ADJ": 37.42, "manlig|ADJ": 37.38, "demonstration|NOUN": 37.37, "färd|NOUN": 37.3, "efterfrågan|NOUN": 37.29, "kandidat|NOUN": 37.23, "upprätthålla|VERB": 37.23, "fördrag|NOUN": 37.17, "instrument|NOUN": 37.17, "analysera|VERB": 37.12, "främmande|ADJ": 37.08, "uppmuntra|VERB": 37.07, "genomförande|NOUN": 37.04, "konservativ|ADJ": 37.03, "attityd|NOUN": 36.99, "föreställning|NOUN": 36.97, "än|SCONJ": 36.96, "lyda|VERB": 36.93, "juridisk|ADJ": 36.89, "variant|NOUN": 36.89, "höjd|NOUN": 36.87, "utrikesminister|NOUN": 36.87, "gäst|NOUN": 36.85, "hustru|NOUN": 36.85, "vandring|NOUN": 36.83, "kontakta|VERB": 36.81, "mil|NOUN": 36.74, "kort|ADV": 36.7, "eventuellt (förk. ev.)|ADV": 36.69, "lära|NOUN": 36.63, "medge|VERB": 36.61, "ologisk|ADJ": 36.6, "alkohol|NOUN": 36.54, "invandring|NOUN": 36.54, "arbetarklass|NOUN": 36.51, "lögn|NOUN": 36.5, "yttrande|NOUN": 36.5, "tillfällig|ADJ": 36.49, "varav|ADV": 36.47, "doktor (förk. dr)|NOUN": 36.39, "olaglig|ADJ": 36.39, "gränsa|VERB": 36.39, "vision|NOUN": 36.38, "framöver|ADV": 36.31, "över|ADV": 36.31, "omgivning|NOUN": 36.28, "bistånd|NOUN": 36.19, "ansluta|VERB": 36.17, "bas|NOUN": 36.17, "fil|NOUN": 36.17, "föredra|VERB": 36.14, "hemma|PART": 36.09, "sönder|PART": 36.03, "etablerad|ADJ": 36.03, "välkomna|VERB": 36.02, "tillverka|VERB": 35.95, "ambition|NOUN": 35.85, "aktie|NOUN": 35.75, "anklaga|VERB": 35.75, "dygn|NOUN": 35.75, "förtjäna|VERB": 35.75, "hur som helst (el. hursomhelst)|ADV": 35.69, "norm|NOUN": 35.69, "osäker|ADJ": 35.63, "räkning|NOUN": 35.61, "republik|NOUN": 35.57, "rykte|NOUN": 35.54, "jämförelse|NOUN": 35.52, "avstå|VERB": 35.46, "ära|NOUN": 35.43, "länsstyrelse|NOUN": 35.41, "smart|ADJ": 35.4, "bibliotek|NOUN": 35.39, "diktatur|NOUN": 35.37, "variera|VERB": 35.35, "dominera|VERB": 35.32, "utreda|VERB": 35.32, "boende|NOUN": 35.29, "museum|NOUN": 35.28, "förvandla|VERB": 35.27, "påbörja|VERB": 35.26, "ursäkt|NOUN": 35.24, "vete|NOUN": 35.23, "organisera|VERB": 35.17, "kommunistisk|ADJ": 35.16, "öra|NOUN": 35.14, "aktivt|ADV": 35.1, "granskning|NOUN": 35.1, "balans|NOUN": 35.09, "mage|NOUN": 35.09, "teckna|VERB": 35.07, "arg|ADJ": 35.03, "säkra|VERB": 35.0, "lunch|NOUN": 34.98, "kommunist|NOUN": 34.92, "militär|NOUN": 34.9, "gåva|NOUN": 34.86, "för närvarande|ADV": 34.84, "alternativ|ADJ": 34.82, "befintlig|ADJ": 34.8, "hälsa|VERB": 34.8, "socialism|NOUN": 34.75, "ursprunglig|ADJ": 34.75, "anställning|NOUN": 34.72, "ansökan|NOUN": 34.66, "protest|NOUN": 34.62, "test|NOUN": 17.8, "anda|NOUN": 34.6, "galen|ADJ": 34.56, "katastrof|NOUN": 34.56, "hata|VERB": 34.52, "gissa|VERB": 34.5, "mur|NOUN": 34.49, "tjänsteman|NOUN": 34.46, "led|NOUN": 8.78, "beakta|VERB": 34.42, "till följd av|ADP": 34.39, "reglera|VERB": 34.32, "kristdemokrat|NOUN": 34.3, "flod|NOUN": 34.29, "talare|NOUN": 34.29, "mörker|NOUN": 34.28, "begränsning|NOUN": 34.27, "värme|NOUN": 34.25, "agerande|NOUN": 34.24, "minoritet|NOUN": 34.2, "etablera|VERB": 34.17, "dam|NOUN": 34.16, "spansk|ADJ": 34.14, "motiv|NOUN": 34.12, "olikhet|NOUN": 34.12, "rättslig|ADJ": 34.11, "utställning|NOUN": 34.11, "utomlands|ADV": 34.1, "huvudstad|NOUN": 34.08, "likt|ADV": 34.08, "terrorist|NOUN": 34.04, "besökare|NOUN": 34.03, "hushåll|NOUN": 34.01, "respektera|VERB": 33.96, "fullständig|ADJ": 33.96, "mäktig|ADJ": 33.88, "växande|ADJ": 33.82, "stabil|ADJ": 33.81, "förvaltning|NOUN": 33.74, "hat|NOUN": 33.72, "mönster|NOUN": 33.72, "nyss|ADV": 33.64, "varumärke|NOUN": 33.62, "fastighet|NOUN": 33.61, "inta|VERB": 33.6, "orolig|ADJ": 33.6, "rulla|VERB": 33.6, "moral|NOUN": 33.59, "motivera|VERB": 33.56, "myt|NOUN": 33.55, "noga|ADV": 33.53, "snacka|VERB": 33.46, "till sist|ADV": 33.46, "förmedla|VERB": 33.45, "hamn|NOUN": 33.39, "tillhandahålla|VERB": 33.37, "informera|VERB": 33.33, "karta|NOUN": 33.33, "utforma|VERB": 33.33, "konvention|NOUN": 33.31, "allt mer (el. alltmer)|ADV": 33.3, "koll|NOUN": 33.3, "längd|NOUN": 33.28, "medicinsk|ADJ": 33.28, "läggning|NOUN": 33.2, "kilogram (el. kilo; förk. kg)|NOUN": 33.17, "finansiering|NOUN": 33.11, "löfte|NOUN": 33.11, "mörda|VERB": 33.11, "anställd|ADJ": 33.1, "amerikan|NOUN": 33.09, "rit|NOUN": 33.09, "status|NOUN": 33.08, "biologisk|ADJ": 33.07, "dikt|NOUN": 33.01, "sko|NOUN": 33.0, "sträcka|VERB": 32.99, "medarbetare|NOUN": 32.96, "lust|NOUN": 32.94, "kassa|NOUN": 32.91, "flygplats|NOUN": 32.9, "tingsrätt|NOUN": 32.89, "avdelning|NOUN": 32.87, "säkerställa|VERB": 32.87, "åklagare|NOUN": 32.84, "lysa|VERB": 32.82, "lidande|NOUN": 32.76, "syna|VERB": 32.75, "standard|NOUN": 32.74, "olycka|NOUN": 32.73, "term|NOUN": 32.71, "maskin|NOUN": 32.7, "transport|NOUN": 32.7, "etisk|ADJ": 32.68, "fattigdom|NOUN": 32.68, "servera|VERB": 32.68, "intern|ADJ": 32.67, "trolig|ADJ": 32.66, "golv|NOUN": 32.64, "förmiddag (förk. fm.)|NOUN": 32.6, "statsråd|NOUN": 32.56, "inrätta|VERB": 32.55, "närhet|NOUN": 32.51, "semester|NOUN": 32.51, "därigenom|ADV": 32.5, "ras|NOUN": 32.4, "tysk|NOUN": 32.38, "favorit|NOUN": 32.27, "framsteg|NOUN": 32.25, "tillvaro|NOUN": 32.25, "faktisk|ADJ": 32.24, "stolt|ADJ": 32.21, "strax|ADV": 32.17, "strida|VERB": 32.17, "angelägen|ADJ": 32.13, "skylla|VERB": 32.1, "ont|ADV": 32.07, "engagera|VERB": 32.0, "beräkning|NOUN": 31.99, "välkommen|ADJ": 31.98, "ideologisk|ADJ": 31.97, "finger|NOUN": 31.96, "hål|NOUN": 31.96, "prövning|NOUN": 31.96, "vettig|ADJ": 31.95, "komplicerad|ADJ": 31.95, "sund|ADJ": 31.91, "domare|NOUN": 31.82, "frukt|NOUN": 31.82, "signal|NOUN": 31.8, "guld|NOUN": 31.79, "homosexuell|ADJ": 31.79, "brottslighet|NOUN": 31.78, "rejäl|ADJ": 31.77, "rättegång|NOUN": 31.75, "mått|NOUN": 31.71, "kammare|NOUN": 31.7, "nazist|NOUN": 31.7, "förefalla|VERB": 31.68, "efteråt|ADV": 31.67, "försäkring|NOUN": 31.67, "konung|NOUN": 31.64, "såklart|ADV": 31.62, "ändamål|NOUN": 31.62, "avsedd|ADJ": 31.62, "generell|ADJ": 31.6, "kommunism|NOUN": 31.6, "dölja|VERB": 31.58, "arab|NOUN": 31.56, "sträva|VERB": 31.5, "stämning|NOUN": 31.5, "torg|NOUN": 31.5, "planerad|ADJ": 31.5, "utrustning|NOUN": 31.48, "vandra|VERB": 31.46, "registrera|VERB": 31.44, "argumentera|VERB": 31.43, "kök|NOUN": 31.43, "uppgå|VERB": 31.41, "visst|INTJ": 31.4, "bön|NOUN": 31.39, "anläggning|NOUN": 31.35, "filosofi|NOUN": 31.35, "gråta|VERB": 31.33, "underlag|NOUN": 31.33, "typisk|ADJ": 31.31, "förespråka|VERB": 31.23, "smärta|NOUN": 31.2, "uppror|NOUN": 31.2, "strategisk|ADJ": 31.17, "symbol|NOUN": 31.17, "radikal|ADJ": 31.16, "VD (verkställande direktör)|NOUN": 31.15, "frid|NOUN": 31.1, "arbetskraft|NOUN": 31.08, "bevilja|VERB": 31.06, "rot|NOUN": 31.06, "förmå|VERB": 31.05, "rak|ADJ": 30.99, "formulera|VERB": 30.98, "jämställdhet|NOUN": 30.98, "existens|NOUN": 30.97, "bonde|NOUN": 30.96, "bränna|VERB": 30.94, "italiensk|ADJ": 30.91, "utgift|NOUN": 30.88, "förbättring|NOUN": 30.87, "föreställa|VERB": 30.83, "operation|NOUN": 30.83, "landa|VERB": 30.82, "service|NOUN": 30.77, "låsa|VERB": 30.76, "varna|VERB": 30.73, "anställa|VERB": 30.69, "förtryck|NOUN": 30.68, "varelse|NOUN": 30.68, "tyst|ADJ": 30.67, "bredvid|ADP": 30.67, "syssla|VERB": 30.67, "drömma|VERB": 30.66, "evangelium|NOUN": 30.61, "planet|NOUN": 30.61, "organiserad|ADJ": 30.6, "fält|NOUN": 30.57, "omröstning|NOUN": 30.56, "psykisk|ADJ": 30.54, "fåtal|NOUN": 30.53, "öppet|ADV": 30.52, "överväga|VERB": 30.52, "stopp|NOUN": 30.49, "tråd|NOUN": 30.46, "prov|NOUN": 30.45, "sinne|NOUN": 30.45, "sorg|NOUN": 30.45, "ensamt|ADV": 30.41, "gemensamt|ADV": 30.41, "bort|ADV": 30.4, "kommersiell|ADJ": 30.4, "före detta (förk. f.d., f d)|ADV": 30.39, "sist|ADV": 30.39, "i huvudsak|ADV": 30.38, "lämpa sig|VERB": 30.37, "annorlunda|ADV": 30.35, "lura|VERB": 30.35, "förvisso|ADV": 30.34, "övervakning|NOUN": 30.33, "pågående|ADJ": 30.32, "utvärdering|NOUN": 30.3, "trygg|ADJ": 30.29, "arv|NOUN": 30.28, "seminarium|NOUN": 30.27, "besvara|VERB": 30.25, "övergrepp|NOUN": 30.21, "pass|NOUN": 30.2, "ljuga|VERB": 30.17, "uppdatering|NOUN": 30.16, "grekisk|ADJ": 30.14, "närvaro|NOUN": 30.09, "tidskrift|NOUN": 30.07, "infrastruktur|NOUN": 30.05, "biskop|NOUN": 30.01, "läger|NOUN": 29.98, "mer och mer|ADV": 29.9, "adress|NOUN": 29.89, "efterhand|ADV": 29.89, "förvånad|ADJ": 29.87, "ovanlig|ADJ": 29.84, "jävla (el. djävla)|ADJ": 29.81, "kontrakt|NOUN": 29.78, "skild|ADJ": 29.77, "daglig|ADJ": 29.75, "penningpolitik|NOUN": 29.75, "röstning|NOUN": 29.75, "lugnt|ADV": 29.74, "video|NOUN": 29.74, "med hänsyn till|ADP": 29.73, "översätta|VERB": 29.68, "fågel|NOUN": 29.62, "inkludera|VERB": 29.6, "era|NOUN": 29.6, "rörande|ADP": 29.57, "förena|VERB": 29.56, "ledig|ADJ": 29.56, "kärnkraft|NOUN": 29.53, "onödig|ADJ": 29.5, "ryss|NOUN": 29.39, "känslig|ADJ": 29.38, "smak|NOUN": 29.35, "order|NOUN": 29.34, "avancerad|ADJ": 29.34, "deltagande|NOUN": 29.32, "nämnd|NOUN": 29.32, "absolut|ADJ": 29.29, "israel|NOUN": 29.29, "prioritera|VERB": 29.23, "tillägga|VERB": 29.23, "blåsa|VERB": 29.2, "trädgård|NOUN": 29.17, "kors|NOUN": 29.16, "nyfiken|ADJ": 29.16, "kombination|NOUN": 29.15, "mod|NOUN": 29.15, "landskap|NOUN": 29.14, "överlämna|VERB": 29.1, "vinnare|NOUN": 29.09, "oskyldig|ADJ": 29.07, "fastna|VERB": 29.01, "förväntning|NOUN": 28.99, "temperatur|NOUN": 28.99, "övergripande|ADJ": 28.98, "motverka|VERB": 28.98, "våldsam|ADJ": 28.97, "fack|NOUN": 28.96, "komplettera|VERB": 28.94, "protokoll|NOUN": 28.94, "webb (el. web)|NOUN": 28.92, "bota|VERB": 28.9, "förlag|NOUN": 28.89, "bege sig|VERB": 28.89, "konsumtion|NOUN": 28.83, "värdefull|ADJ": 28.83, "kost|NOUN": 28.82, "godkänd|ADJ": 28.82, "datum|NOUN": 28.69, "därtill|ADV": 28.65, "recension|NOUN": 28.65, "till|ADV": 28.65, "omsorg|NOUN": 28.61, "kriterium|NOUN": 28.6, "fånge|NOUN": 28.6, "extrem|ADJ": 28.56, "förbindelse|NOUN": 28.54, "angrepp|NOUN": 28.53, "lansera|VERB": 28.52, "saga|NOUN": 28.5, "basera|VERB": 28.48, "cykel|NOUN": 28.46, "design|NOUN": 28.45, "frivillig|ADJ": 28.45, "med anledning av|ADP": 28.44, "västra|ADJ": 28.43, "påverkan|NOUN": 28.4, "verkan|NOUN": 28.4, "ful|ADJ": 28.39, "kongress|NOUN": 28.37, "skära|VERB": 28.35, "testamente|NOUN": 28.35, "gul|ADJ": 28.34, "skriftlig|ADJ": 28.34, "våg|NOUN": 28.31, "årlig|ADJ": 28.31, "reservation|NOUN": 28.25, "rättvis|ADJ": 28.24, "yrke|NOUN": 28.24, "århundrade|NOUN": 28.24, "anslag|NOUN": 28.22, "drog|NOUN": 28.17, "gömma|VERB": 28.13, "äkta|ADJ": 28.13, "intellektuell|ADJ": 28.09, "kejsare|NOUN": 28.05, "planering|NOUN": 28.05, "släkt|NOUN": 27.98, "drottning|NOUN": 27.97, "uppträda|VERB": 27.94, "övergå|VERB": 27.94, "het|ADJ": 27.88, "läkemedel|NOUN": 27.87, "utformning|NOUN": 27.85, "elektronisk|ADJ": 27.83, "obligatorisk|ADJ": 27.76, "investera|VERB": 27.72, "fond|NOUN": 27.71, "dubbel|ADJ": 27.69, "uppkomma|VERB": 27.67, "somna|VERB": 27.63, "ställningstagande|NOUN": 27.63, "utesluta|VERB": 27.6, "frukost|NOUN": 27.59, "förhoppning|NOUN": 27.59, "facklig|ADJ": 27.56, "prognos|NOUN": 27.55, "sannolikhet|NOUN": 27.54, "advokat|NOUN": 27.53, "kapitalistisk|ADJ": 27.52, "tveksam|ADJ": 27.46, "anlända|VERB": 27.46, "regn|NOUN": 27.44, "röja|VERB": 27.4, "motsats|NOUN": 27.39, "referens|NOUN": 27.39, "fabrik|NOUN": 27.37, "i och för sig|ADV": 27.37, "japansk|ADJ": 27.32, "plus|ADV": 27.31, "marknadsföring|NOUN": 27.3, "rena|VERB": 27.3, "innebörd|NOUN": 27.24, "stjäla|VERB": 27.23, "online|ADV": 27.21, "omgång|NOUN": 27.19, "protestera|VERB": 27.17, "tillkomma|VERB": 27.17, "bemöta|VERB": 27.15, "tränga|VERB": 27.15, "bestående|ADJ": 27.11, "blomma|NOUN": 27.1, "överföra|VERB": 27.1, "solidaritet|NOUN": 27.1, "lydelse|NOUN": 27.08, "annons|NOUN": 27.05, "riksdagsledamot|NOUN": 27.04, "brinna|VERB": 27.03, "rinna|VERB": 27.03, "gärning|NOUN": 27.03, "samverkan|NOUN": 27.03, "rymma|VERB": 27.01, "blogginlägg|NOUN": 27.0, "sammanfatta|VERB": 26.98, "östra|ADJ": 26.97, "dröja|VERB": 26.96, "avbryta|VERB": 26.95, "gräva|VERB": 26.93, "stryka|VERB": 26.93, "kreativ|ADJ": 26.92, "till dess|ADV": 26.91, "intensiv|ADJ": 26.9, "sålunda|ADV": 26.84, "roa|VERB": 26.83, "understryka|VERB": 26.82, "glas|NOUN": 26.81, "album|NOUN": 26.79, "territorium|NOUN": 26.78, "möjliggöra|VERB": 26.75, "fördelning|NOUN": 26.74, "folkomröstning|NOUN": 26.74, "skede|NOUN": 26.73, "markera|VERB": 26.72, "skaka|VERB": 26.71, "sten|NOUN": 26.71, "vagn|NOUN": 26.71, "värna|VERB": 26.7, "hemsk|ADJ": 26.68, "kriminell|ADJ": 26.67, "saklig|ADJ": 26.64, "närvarande|ADJ": 26.63, "automatiskt|ADV": 26.61, "skämma|VERB": 26.61, "vittna|VERB": 26.6, "spendera|VERB": 26.6, "ansvara|VERB": 26.59, "ledarskap|NOUN": 26.59, "trivas|VERB": 26.58, "figur|NOUN": 26.57, "bygd|NOUN": 26.56, "spridning|NOUN": 26.56, "lyckad|ADJ": 26.55, "le|VERB": 26.54, "betalning|NOUN": 26.52, "oroa|VERB": 26.52, "lov|NOUN": 26.46, "motsatt|ADJ": 26.46, "knyta|VERB": 26.45, "från och med|ADP": 26.44, "rekommendation|NOUN": 26.44, "ansträngning|NOUN": 26.41, "institut|NOUN": 26.41, "kritiker|NOUN": 26.41, "övre|ADJ": 26.39, "moderat|ADJ": 26.38, "data|NOUN": 26.32, "hörn|NOUN": 26.31, "inhemsk|ADJ": 26.31, "öl|NOUN": 26.31, "ängel|NOUN": 26.29, "blott|ADV": 26.28, "förhålla sig|VERB": 26.27, "förhålla|VERB": 26.27, "park|NOUN": 26.25, "regelverk|NOUN": 26.23, "nackdel|NOUN": 26.22, "vittne|NOUN": 26.21, "ljus|ADJ": 26.17, "medvetet|ADV": 26.15, "gas|NOUN": 26.13, "tipsa|VERB": 26.13, "våldtäkt|NOUN": 26.11, "boka|VERB": 26.1, "sådan här (vardagl. sån här)|DET": 26.09, "ekologisk|ADJ": 26.08, "återfinna|VERB": 26.08, "huvudsakligen|ADV": 26.07, "överge|VERB": 26.04, "ockupation|NOUN": 26.03, "likaså|ADV": 26.02, "bringa|VERB": 26.0, "hylla|VERB": 25.98, "sammanfattning|NOUN": 25.98, "liberal|NOUN": 25.97, "graf|NOUN": 25.96, "slott|NOUN": 25.96, "anspråk|NOUN": 25.94, "motsättning|NOUN": 25.92, "byte|NOUN": 25.89, "logik|NOUN": 25.88, "resonera|VERB": 25.87, "tempel|NOUN": 25.85, "krönika|NOUN": 25.84, "tillbringa|VERB": 25.83, "kopia|NOUN": 25.82, "instans|NOUN": 25.8, "företagare|NOUN": 25.78, "medlemskap|NOUN": 25.76, "egentlig|ADJ": 25.75, "landsbygd|NOUN": 25.75, "integration|NOUN": 25.74, "gest|NOUN": 25.74, "tyst|ADV": 25.74, "längta|VERB": 25.72, "föreskrift|NOUN": 25.67, "generellt|ADV": 25.67, "konto|NOUN": 25.67, "ju|CCONJ": 25.65, "tämligen|ADV": 25.65, "då och då|ADV": 25.64, "ryka|VERB": 25.61, "reglering|NOUN": 25.6, "misstänkt|ADJ": 25.55, "paket|NOUN": 25.51, "bete sig|VERB": 25.49, "kollektiv|ADJ": 25.48, "fotograf|NOUN": 25.47, "vänlig|ADJ": 25.46, "hemlighet|NOUN": 25.45, "administrativ|ADJ": 25.42, "dansa|VERB": 25.41, "tillägg|NOUN": 25.41, "fordon|NOUN": 25.4, "nöja sig|VERB": 25.39, "kliva|VERB": 25.38, "bro|NOUN": 25.37, "mandat|NOUN": 25.35, "inledning|NOUN": 25.34, "införande|NOUN": 25.33, "antyda|VERB": 25.32, "innefatta|VERB": 25.32, "kommunicera|VERB": 25.32, "praktiskt|ADV": 25.32, "förmån|NOUN": 25.31, "motivering|NOUN": 25.31, "tystnad|NOUN": 25.3, "valuta|NOUN": 25.29, "genomgå|VERB": 25.25, "nåd|NOUN": 25.24, "redaktion|NOUN": 25.24, "extern|ADJ": 25.22, "sfär|NOUN": 25.22, "flygplan|NOUN": 25.2, "kamrat|NOUN": 25.18, "premiärminister|NOUN": 25.18, "botten|NOUN": 25.17, "västerländsk|ADJ": 25.17, "skala|NOUN": 25.14, "utsikt|NOUN": 25.14, "besegra|VERB": 25.12, "utfärda|VERB": 25.12, "stimulera|VERB": 25.1, "kraftfull|ADJ": 25.03, "utöka|VERB": 25.03, "angripa|VERB": 25.02, "utseende|NOUN": 25.02, "promenad|NOUN": 25.0, "universum|NOUN": 24.97, "vanligtvis|ADV": 24.95, "pensionär|NOUN": 24.91, "redo|ADJ": 24.9, "järnväg|NOUN": 24.89, "jämn|ADJ": 24.89, "utbyte|NOUN": 24.89, "öppenhet|NOUN": 24.89, "grundval|NOUN": 24.88, "attackera|VERB": 24.87, "slita|VERB": 24.84, "förskola|NOUN": 24.83, "föregående|ADJ": 24.82, "föreskriva|VERB": 24.82, "inspiration|NOUN": 24.82, "anhängare|NOUN": 24.82, "hyra|VERB": 24.8, "kärna|NOUN": 24.79, "över huvud taget (el. överhuvudtaget)|ADV": 24.79, "löpa|VERB": 24.75, "blad|NOUN": 24.74, "gårdag|NOUN": 24.73, "tillföra|VERB": 24.71, "trovärdighet|NOUN": 24.71, "varv|NOUN": 24.71, "värdighet|NOUN": 24.71, "dans|NOUN": 24.7, "osäkerhet|NOUN": 24.7, "enstaka|ADJ": 24.69, "flyg|NOUN": 24.66, "vana|NOUN": 24.66, "spänning|NOUN": 24.64, "anfall|NOUN": 24.63, "utarbeta|VERB": 24.62, "skrämma|VERB": 24.6, "nyckel|NOUN": 24.59, "skribent|NOUN": 24.54, "garanti|NOUN": 24.53, "sakta|ADV": 24.53, "tillsätta|VERB": 24.51, "tvekan|NOUN": 24.51, "tand|NOUN": 24.5, "yrka|VERB": 24.5, "tacksam|ADJ": 24.47, "tävla|VERB": 24.44, "bortom|ADP": 24.39, "utbilda|VERB": 24.39, "hemland|NOUN": 24.39, "utav|ADP": 24.37, "avvisa|VERB": 24.36, "potentiell|ADJ": 24.32, "sovjetisk|ADJ": 24.3, "skepp|NOUN": 24.29, "utgång|NOUN": 24.25, "skrämmande|ADJ": 24.23, "omedelbar|ADJ": 24.21, "partner|NOUN": 24.16, "rejält|ADV": 24.12, "kapacitet|NOUN": 24.06, "genomsnitt|NOUN": 24.04, "värdig|ADJ": 24.02, "gymnasium|NOUN": 24.0, "umgås|VERB": 23.99, "knä|NOUN": 23.97, "element|NOUN": 23.96, "fredlig|ADJ": 23.96, "smal|ADJ": 23.96, "gubbe|NOUN": 23.96, "arrangera|VERB": 23.95, "skugga|NOUN": 23.95, "pressa|VERB": 23.86, "självständighet|NOUN": 23.85, "densamma|PRON": 23.84, "slutlig|ADJ": 23.83, "tvivel|NOUN": 23.82, "fälla|VERB": 23.8, "smaka|VERB": 23.78, "näst|ADV": 23.75, "utbud|NOUN": 23.75, "opinion|NOUN": 23.75, "värdera|VERB": 23.75, "allvarligt|ADV": 23.74, "formell|ADJ": 23.74, "dagligen|ADV": 23.71, "ursprungligen|ADV": 23.71, "vidare|ADJ": 23.71, "fördela|VERB": 23.67, "ovanligt|ADV": 23.67, "reducera|VERB": 23.67, "vanligt|ADV": 23.67, "skadestånd|NOUN": 23.63, "kopiera|VERB": 23.62, "övergång|NOUN": 23.6, "anhörig|ADJ": 23.6, "ångest|NOUN": 23.6, "vakt|NOUN": 23.59, "förhandla|VERB": 23.58, "koncentrera|VERB": 23.58, "tabell|NOUN": 23.57, "önskan|NOUN": 23.53, "konsert|NOUN": 23.52, "teckning|NOUN": 23.51, "avgå|VERB": 23.46, "grav|NOUN": 23.45, "agenda|NOUN": 23.43, "samfund|NOUN": 23.4, "krets|NOUN": 23.39, "kunglig|ADJ": 23.37, "anmälan|NOUN": 23.34, "inneha|VERB": 23.34, "soffa|NOUN": 23.32, "stabilitet|NOUN": 23.32, "förnuft|NOUN": 23.3, "därav|ADV": 23.28, "tredjedel|NOUN": 23.27, "ovanstående|ADJ": 23.26, "trovärdig|ADJ": 23.26, "strunta|VERB": 23.24, "akademisk|ADJ": 23.23, "permanent|ADJ": 23.23, "nyttig|ADJ": 23.2, "invändning|NOUN": 23.17, "våning|NOUN": 23.11, "långsamt|ADV": 23.1, "vild|ADJ": 23.1, "propaganda|NOUN": 23.09, "troende|ADJ": 23.07, "exemplar|NOUN": 23.05, "resolution|NOUN": 23.04, "ekonomiskt|ADV": 23.03, "därpå|ADV": 23.03, "formulering|NOUN": 23.03, "ihjäl|PART": 23.01, "såväl som|CCONJ": 23.0, "instämma|VERB": 22.98, "halvår|NOUN": 22.97, "debattera|VERB": 22.96, "idiot|NOUN": 22.96, "yttersta|ADJ": 22.96, "intill|ADP": 22.95, "torr|ADJ": 22.93, "söt|ADJ": 22.92, "socialist|NOUN": 22.91, "anordna|VERB": 22.9, "besviken|ADJ": 22.89, "lektion|NOUN": 22.89, "ledsen|ADJ": 22.86, "grattis|INTJ": 22.84, "sistnämnd|ADJ": 22.83, "tragisk|ADJ": 22.83, "teater|NOUN": 22.82, "försäkra|VERB": 22.81, "ideal|NOUN": 22.81, "vice|ADJ": 22.81, "hantering|NOUN": 22.8, "målsättning|NOUN": 22.78, "begripa|VERB": 22.77, "upphov|NOUN": 22.74, "kränka|VERB": 22.72, "i morse (el. imorse)|ADV": 22.71, "hals|NOUN": 22.7, "mån|NOUN": 22.7, "stam|NOUN": 22.7, "journalistik|NOUN": 22.67, "intäkt|NOUN": 22.66, "mjuk|ADJ": 22.66, "Bproper name (bruttonationalprodukt)|NOUN": 22.63, "grå|ADJ": 22.63, "profil|NOUN": 22.61, "krossa|VERB": 22.6, "partiledare|NOUN": 22.6, "centimeter (förk. cm)|NOUN": 22.59, "övertyga|VERB": 22.59, "romersk|ADJ": 22.56, "sörja|VERB": 22.56, "inspirera|VERB": 22.55, "övertygelse|NOUN": 22.54, "stackars|ADJ": 22.52, "sänkning|NOUN": 22.5, "potential|NOUN": 22.48, "antagande|NOUN": 22.47, "tilldela|VERB": 22.46, "biljett|NOUN": 22.43, "motsätta|VERB": 22.41, "komplex|ADJ": 22.4, "skadad|ADJ": 22.39, "begäran|NOUN": 22.38, "arena|NOUN": 22.36, "kust|NOUN": 22.36, "åtal|NOUN": 22.36, "dimension|NOUN": 22.34, "internationellt|ADV": 22.34, "nationellt|ADV": 22.34, "hållning|NOUN": 22.33, "gen|NOUN": 22.32, "lugn|NOUN": 22.32, "döpa|VERB": 22.32, "fantasi|NOUN": 22.32, "spets|NOUN": 22.3, "avsätta|VERB": 22.29, "fundering|NOUN": 22.29, "kombinera|VERB": 22.27, "observera|VERB": 22.24, "intressera|VERB": 22.23, "uppåt|ADV": 22.23, "fas|NOUN": 22.22, "dop|NOUN": 22.21, "professionell|ADJ": 22.2, "klippa|VERB": 22.18, "trist|ADJ": 22.17, "ombord|ADV": 22.17, "sparka|VERB": 22.17, "klimatförändring|NOUN": 22.16, "undervisa|VERB": 22.14, "dåvarande|ADJ": 22.13, "varning|NOUN": 22.13, "ton|NOUN": 14.81, "tänkbar|ADJ": 22.11, "villig|ADJ": 22.1, "station|NOUN": 22.08, "släkting|NOUN": 22.07, "övrigt|ADV": 22.04, "giltig|ADJ": 22.03, "gudomlig|ADJ": 22.02, "objektiv|ADJ": 22.0, "brand|NOUN": 21.99, "meningslös|ADJ": 21.89, "yttra|VERB": 21.89, "minskning|NOUN": 21.87, "axel|NOUN": 21.84, "försämra|VERB": 21.83, "motor|NOUN": 21.82, "i och med|ADV": 21.81, "konstruktion|NOUN": 21.81, "arkiv|NOUN": 21.8, "äventyr|NOUN": 21.8, "oj|INTJ": 21.78, "Sverige|PROPN": 21.76, "humor|NOUN": 21.75, "like|NOUN": 21.73, "paragraf|NOUN": 21.73, "odla|VERB": 21.69, "erbjudande|NOUN": 21.68, "vidga|VERB": 21.68, "volym|NOUN": 21.67, "motsätta sig|VERB": 21.67, "missbruk|NOUN": 21.66, "utvidga|VERB": 21.64, "snarast|ADV": 21.6, "uppmaning|NOUN": 21.58, "kram|NOUN": 21.56, "intervjua|VERB": 21.55, "livsmedel|NOUN": 21.55, "anklagelse|NOUN": 21.54, "cykla|VERB": 21.54, "samordning|NOUN": 21.54, "dessvärre|ADV": 21.51, "oklar|ADJ": 21.51, "företeelse|NOUN": 21.46, "offra|VERB": 21.46, "lager|NOUN": 21.45, "arbetsliv|NOUN": 21.44, "lysande|ADJ": 21.43, "bränsle|NOUN": 21.4, "finanskris|NOUN": 21.4, "nödvändigtvis|ADV": 21.4, "gott om|ADV": 21.39, "medeltid|NOUN": 21.39, "strävan|NOUN": 21.39, "hastighet|NOUN": 21.38, "kö|NOUN": 21.38, "medvetande|NOUN": 21.37, "producent|NOUN": 21.37, "så pass|ADV": 21.37, "vetande|NOUN": 21.37, "i mitten av|ADP": 21.36, "dylik|ADJ": 21.33, "installera|VERB": 21.32, "utge|VERB": 21.3, "förberedelse|NOUN": 21.28, "fördom|NOUN": 21.25, "synnerligen|ADV": 21.25, "i närheten av|ADP": 21.22, "åtagande|NOUN": 21.22, "tillkännage|VERB": 21.2, "kaos|NOUN": 21.17, "mästare|NOUN": 21.16, "utmana|VERB": 21.16, "drift|NOUN": 21.15, "hundratal|NOUN": 21.15, "måne|NOUN": 21.13, "bita|VERB": 21.11, "blandad|ADJ": 21.1, "hjälte|NOUN": 21.1, "skänka|VERB": 21.09, "tillämplig|ADJ": 21.09, "betydelsefull|ADJ": 21.08, "synsätt|NOUN": 21.07, "ström|NOUN": 21.03, "förse|VERB": 21.02, "mätning|NOUN": 21.02, "massiv|ADJ": 21.01, "atmosfär|NOUN": 20.97, "mall|NOUN": 20.96, "personlighet|NOUN": 20.96, "gren|NOUN": 20.95, "väldig|ADJ": 20.93, "effektivt|ADV": 20.89, "vanligen|ADV": 20.88, "koncept|NOUN": 20.85, "välkänd|ADJ": 20.84, "förebild|NOUN": 20.81, "uppenbart|ADV": 20.81, "recept|NOUN": 20.79, "föreläsning|NOUN": 20.77, "antisemitism|NOUN": 20.75, "geografisk|ADJ": 20.75, "grafisk|ADJ": 20.75, "upplysning|NOUN": 20.74, "general|NOUN": 20.73, "administration|NOUN": 20.72, "bröst|NOUN": 20.69, "tills|ADP": 20.69, "patent|NOUN": 20.67, "befogenhet|NOUN": 20.67, "skarp|ADJ": 20.63, "islamisk|ADJ": 20.6, "vem som helst|PRON": 20.6, "förverkliga|VERB": 20.57, "prioritering|NOUN": 20.57, "vistas|VERB": 20.55, "regelbundet|ADV": 20.53, "depression|NOUN": 20.49, "effektivitet|NOUN": 20.48, "inne|PART": 20.48, "likväl|ADV": 20.48, "blandning|NOUN": 20.47, "datera|VERB": 20.46, "final|NOUN": 20.45, "tjock|ADJ": 20.45, "erövra|VERB": 20.43, "höger|NOUN": 20.43, "sträcka|NOUN": 20.42, "vaka|VERB": 20.41, "polsk|ADJ": 20.4, "bomb|NOUN": 20.39, "tår|NOUN": 20.39, "fackförening|NOUN": 20.37, "utvald|ADJ": 20.36, "placering|NOUN": 20.32, "huvudsaklig|ADJ": 20.31, "avfall|NOUN": 20.3, "gigantisk|ADJ": 20.3, "väntan|NOUN": 20.3, "turnering|NOUN": 20.28, "uppvärmning|NOUN": 20.28, "djup|NOUN": 20.27, "praxis|NOUN": 20.26, "okej|INTJ": 20.25, "maximal (förk. max.)|ADJ": 20.23, "konstitution|NOUN": 20.22, "otrolig|ADJ": 20.22, "fruktansvärd|ADJ": 20.21, "straffa|VERB": 20.2, "sådär|ADV": 20.2, "nödvändighet|NOUN": 20.18, "medlemsland|NOUN": 20.17, "översyn|NOUN": 20.16, "blind|ADJ": 20.15, "front|NOUN": 20.15, "fördöma|VERB": 20.13, "synlig|ADJ": 20.12, "fint|ADV": 20.11, "skapelse|NOUN": 20.1, "rasa|VERB": 20.1, "verksam|ADJ": 20.1, "avlida|VERB": 20.09, "fullkomligt|ADV": 20.09, "teoretisk|ADJ": 20.09, "flyta|VERB": 20.08, "urval|NOUN": 20.07, "binda|VERB": 20.05, "fett|NOUN": 20.03, "erkännande|NOUN": 20.03, "hälsning|NOUN": 20.03, "idrott|NOUN": 20.03, "debattartikel|NOUN": 20.02, "belysa|VERB": 20.0, "emellan|ADP": 19.99, "övervaka|VERB": 19.98, "lagom|ADV": 19.96, "sömn|NOUN": 19.96, "proletariat|NOUN": 19.91, "önskemål|NOUN": 19.91, "förlåta|VERB": 19.89, "sammanlagt|ADV": 19.89, "slav|NOUN": 19.89, "näsa|NOUN": 19.88, "däribland|ADV": 19.85, "export|NOUN": 19.85, "nedgång|NOUN": 19.83, "vinkel|NOUN": 19.83, "experiment|NOUN": 19.82, "allierad|ADJ": 19.81, "arbetstid|NOUN": 19.81, "flagga|NOUN": 19.81, "uppdatera|VERB": 19.81, "block|NOUN": 19.79, "feminism|NOUN": 19.78, "skattebetalare|NOUN": 19.78, "globalisering|NOUN": 19.77, "miljontals|ADV": 19.77, "obehaglig|ADJ": 19.77, "ondska|NOUN": 19.75, "önskvärd|ADJ": 19.74, "anpassad|ADJ": 19.74, "mysig|ADJ": 19.7, "norr|NOUN": 19.7, "andning|NOUN": 19.68, "motta|VERB": 19.68, "utspela sig|VERB": 19.66, "exakt|ADJ": 19.65, "elit|NOUN": 19.64, "inverkan|NOUN": 19.64, "akut|ADJ": 19.61, "kvarstå|VERB": 19.61, "troligtvis|ADV": 19.6, "konkurs|NOUN": 19.58, "center|NOUN": 19.56, "än så länge|ADV": 19.56, "dramatisk|ADJ": 19.55, "låtsas|VERB": 19.54, "underlig|ADJ": 19.54, "förlängning|NOUN": 19.52, "segla|VERB": 19.51, "försiktig|ADJ": 19.5, "himla|ADV": 19.5, "inbördeskrig|NOUN": 19.48, "vid sidan av|ADP": 19.48, "grym|ADJ": 19.47, "tunn|ADJ": 19.47, "grundlag|NOUN": 19.46, "realistisk|ADJ": 19.45, "tvätta|VERB": 19.45, "enormt|ADV": 19.42, "litterär|ADJ": 19.42, "mobiltelefon|NOUN": 19.41, "dominerande|ADJ": 19.38, "framkomma|VERB": 19.38, "misshandel|NOUN": 19.37, "skildra|VERB": 19.34, "förbannad|ADJ": 19.34, "anpassning|NOUN": 19.33, "redaktör|NOUN": 19.31, "behörig|ADJ": 19.3, "last|NOUN": 19.29, "arbetarrörelse|NOUN": 19.28, "liberalism|NOUN": 19.28, "presentation|NOUN": 19.28, "stress|NOUN": 19.27, "försörja|VERB": 19.26, "objekt|NOUN": 19.26, "omslag|NOUN": 19.25, "absurd|ADJ": 19.24, "kvalificerad|ADJ": 19.24, "trappa|NOUN": 19.22, "offentligt|ADV": 19.2, "röka|VERB": 19.2, "valrörelse|NOUN": 19.2, "anfalla|VERB": 19.19, "rådande|ADJ": 19.17, "spåra|VERB": 19.17, "upplaga|NOUN": 19.17, "ordentlig|ADJ": 19.16, "klä (el. kläda)|VERB": 19.15, "ambassad|NOUN": 19.1, "konkurrera|VERB": 19.1, "ovanför|ADP": 19.1, "skämt|NOUN": 19.1, "tända|VERB": 19.1, "anslutning|NOUN": 19.09, "backa|VERB": 19.09, "loss|PART": 19.06, "samvete|NOUN": 19.05, "fastän|SCONJ": 19.04, "årtionde|NOUN": 19.04, "tomt|NOUN": 19.02, "avsevärt|ADV": 19.01, "rita|VERB": 19.01, "värt|ADV": 19.01, "register|NOUN": 19.0, "rörlighet|NOUN": 19.0, "ignorera|VERB": 18.99, "dold|ADJ": 18.98, "befria|VERB": 18.98, "först och främst|ADV": 18.98, "retorik|NOUN": 18.97, "leende|NOUN": 18.95, "olycklig|ADJ": 18.92, "säkerligen|ADV": 18.92, "abort|NOUN": 18.89, "taktik|NOUN": 18.89, "beteckna|VERB": 18.88, "lärjunge|NOUN": 18.88, "stadga|NOUN": 18.87, "långsam|ADJ": 18.86, "oberoende av|ADP": 18.86, "utlänning|NOUN": 18.84, "spelning|NOUN": 18.82, "godkännande|NOUN": 18.8, "fet|ADJ": 18.78, "hovrätt|NOUN": 18.78, "tiotal|NOUN": 18.77, "skivbolag|NOUN": 18.75, "stycke|NOUN": 18.73, "tempo|NOUN": 18.73, "påve|NOUN": 18.7, "kant|NOUN": 18.68, "turist|NOUN": 18.67, "predika|VERB": 18.66, "reflektera|VERB": 18.65, "folkgrupp|NOUN": 18.63, "rektor|NOUN": 18.62, "klargöra|VERB": 18.6, "neutral|ADJ": 18.6, "laglig|ADJ": 18.6, "tendera|VERB": 18.6, "utrikespolitik|NOUN": 18.6, "glädja|VERB": 18.59, "rödgrön|ADJ": 18.56, "segra|VERB": 18.55, "inrikta|VERB": 18.53, "monopol|NOUN": 18.53, "konkurrent|NOUN": 18.52, "plattform|NOUN": 18.51, "skådespelare|NOUN": 18.51, "störning|NOUN": 18.5, "remissinstans|NOUN": 18.47, "rutin|NOUN": 18.47, "dal|NOUN": 18.46, "studio|NOUN": 18.46, "användbar|ADJ": 18.45, "lagförslag|NOUN": 18.45, "självfallet|ADV": 18.45, "ömsesidig|ADJ": 18.43, "förvåna|VERB": 18.41, "flaska|NOUN": 18.39, "packa|VERB": 18.38, "reportage|NOUN": 18.34, "skylt|NOUN": 18.33, "platta|NOUN": 18.32, "välsignelse|NOUN": 18.32, "cell|NOUN": 18.3, "i förväg|ADV": 18.28, "kopp|NOUN": 18.26, "bortse|VERB": 18.25, "etik|NOUN": 18.25, "mördare|NOUN": 18.25, "med stöd av|ADP": 18.24, "vid|ADJ": 18.24, "förintelse|NOUN": 18.23, "redogöra|VERB": 18.23, "auktoritet|NOUN": 18.22, "avslå|VERB": 18.22, "hud|NOUN": 18.22, "välstånd|NOUN": 18.21, "rättfärdig|ADJ": 18.2, "därvid|ADV": 18.19, "tillgodose|VERB": 18.19, "mental|ADJ": 18.19, "försvarsmakt|NOUN": 18.17, "kollektivavtal|NOUN": 18.16, "svaghet|NOUN": 18.16, "frågeställning|NOUN": 18.15, "motsvarighet|NOUN": 18.14, "slutändan|NOUN": 18.14, "bitter|ADJ": 18.13, "utanförskap|NOUN": 18.13, "åtskillig|ADJ": 18.1, "koldioxid|NOUN": 18.08, "mässa|NOUN": 18.08, "rå|ADJ": 18.07, "tvivla|VERB": 18.06, "höjning|NOUN": 18.05, "forn|ADJ": 18.04, "konjunktur|NOUN": 18.03, "nöje|NOUN": 18.03, "attraktiv|ADJ": 17.99, "reflektion|NOUN": 17.99, "samråd|NOUN": 17.97, "afrikansk|ADJ": 17.96, "kontroversiell|ADJ": 17.96, "ruta|NOUN": 17.96, "folklig|ADJ": 17.94, "framträda|VERB": 17.93, "vis|ADJ": 17.93, "förlänga|VERB": 17.92, "spegla|VERB": 17.91, "frånvaro|NOUN": 17.9, "symptom (el. symtom)|NOUN": 17.9, "bokstav|NOUN": 17.89, "webbläsare|NOUN": 17.85, "skrivelse|NOUN": 17.84, "barndom|NOUN": 17.83, "usel|ADJ": 17.81, "folkmord|NOUN": 17.8, "till känna|ADV": 17.8, "arbetsuppgift|NOUN": 17.78, "illegal|ADJ": 17.78, "städa|VERB": 17.78, "uppvisa|VERB": 17.78, "väska|NOUN": 17.78, "ärligt|ADV": 17.78, "historiskt|ADV": 17.76, "upphovsman|NOUN": 17.76, "lock|NOUN": 17.75, "tes|NOUN": 17.75, "bekostnad|NOUN": 17.74, "info|NOUN": 17.74, "skadlig|ADJ": 17.74, "ansöka|VERB": 17.73, "industriell|ADJ": 17.73, "köpare|NOUN": 17.73, "börs|NOUN": 17.72, "beklaga|VERB": 17.7, "korruption|NOUN": 17.66, "uppföra|VERB": 17.66, "arbetsförmedling|NOUN": 17.65, "fria|VERB": 17.65, "britt|NOUN": 17.64, "kontinent|NOUN": 17.64, "låda|NOUN": 17.64, "bevaka|VERB": 17.61, "besparing|NOUN": 17.6, "redovisning|NOUN": 17.59, "variation|NOUN": 17.59, "detaljerad|ADJ": 17.59, "skratt|NOUN": 17.58, "naken|ADJ": 17.56, "byggande|NOUN": 17.54, "konstruktiv|ADJ": 17.53, "integrera|VERB": 17.5, "återkommande|ADJ": 17.49, "slump|NOUN": 17.49, "mottagare|NOUN": 17.47, "återgå|VERB": 17.47, "i likhet med|ADV": 17.46, "leverantör|NOUN": 17.46, "noll|NUM": 17.45, "storm|NOUN": 17.45, "pirat|NOUN": 17.42, "svänga|VERB": 17.42, "bifall|NOUN": 17.41, "instruktion|NOUN": 17.39, "upptagen|ADJ": 17.39, "paus|NOUN": 17.37, "rationell|ADJ": 17.36, "överstiga|VERB": 17.36, "delad|ADJ": 17.35, "skärpa|VERB": 17.35, "tillverkare|NOUN": 17.34, "imponerande|ADJ": 17.34, "följaktligen|ADV": 17.32, "innan|ADP": 17.32, "misstanke|NOUN": 17.32, "omdöme|NOUN": 17.32, "kod|NOUN": 17.31, "server|NOUN": 17.31, "magisk|ADJ": 17.29, "sträng|ADJ": 17.29, "vad som helst|ADV": 17.27, "dagbok|NOUN": 17.25, "radera|VERB": 17.25, "anknytning|NOUN": 17.23, "häromdagen|ADV": 17.23, "innovation|NOUN": 17.23, "gran|NOUN": 17.21, "uppföljning|NOUN": 17.21, "grabb|NOUN": 17.2, "frukta|VERB": 17.18, "tvist|NOUN": 17.16, "innan|ADV": 17.15, "van|ADJ": 17.15, "dubbelt|ADV": 17.14, "mild|ADJ": 17.14, "drivkraft|NOUN": 17.11, "tjänare|NOUN": 17.09, "nationalism|NOUN": 17.08, "moln|NOUN": 17.07, "ordförandeskap|NOUN": 17.07, "såvitt|SCONJ": 17.07, "mekanism|NOUN": 17.06, "minsann|ADV": 17.06, "vaccin|NOUN": 17.06, "filosof|NOUN": 17.05, "division|NOUN": 17.03, "belägen|ADJ": 17.02, "tåla|VERB": 17.01, "avdrag|NOUN": 17.0, "koloni|NOUN": 17.0, "sannerligen|ADV": 17.0, "till förmån för|ADP": 16.96, "cancer|NOUN": 16.95, "förföljelse|NOUN": 16.95, "byråkrati|NOUN": 16.94, "mobil|ADJ": 16.93, "tillsyn|NOUN": 16.93, "ett|PRON": 16.92, "sur|ADJ": 16.92, "nazism|NOUN": 16.9, "rösträtt|NOUN": 16.89, "somlig|PRON": 16.89, "utredare|NOUN": 16.89, "stadium|NOUN": 16.88, "dagis|NOUN": 16.87, "färsk|ADJ": 16.86, "positivt|ADV": 16.86, "livsstil|NOUN": 16.85, "pressmeddelande|NOUN": 16.83, "klyfta|NOUN": 16.82, "skapande|NOUN": 16.82, "inlagd|ADJ": 16.82, "konstnärlig|ADJ": 16.81, "pinsam|ADJ": 16.81, "löpande|ADJ": 16.8, "konstant|ADJ": 16.8, "åberopa|VERB": 16.8, "arrangemang|NOUN": 16.78, "avslutad|ADJ": 16.78, "varifrån|ADV": 16.77, "jurist|NOUN": 16.76, "lagra|VERB": 16.75, "påtaglig|ADJ": 16.75, "tillgänglighet|NOUN": 16.75, "pedagogisk|ADJ": 16.73, "skita|VERB": 16.73, "kärnvapen|NOUN": 16.71, "plikt|NOUN": 16.71, "företräda|VERB": 16.68, "mjölk|NOUN": 16.68, "policy|NOUN": 16.68, "ångra|VERB": 16.66, "apostel|NOUN": 16.65, "ingripa|VERB": 16.64, "tröttna|VERB": 16.63, "utvidgning|NOUN": 16.63, "kvarter|NOUN": 16.62, "flexibel|ADJ": 16.61, "motionär|NOUN": 16.6, "ideell|ADJ": 16.58, "insyn|NOUN": 16.58, "bosatt|ADJ": 16.57, "filosofisk|ADJ": 16.54, "inspelning|NOUN": 16.53, "reell|ADJ": 16.53, "generera|VERB": 16.53, "krypa|VERB": 16.5, "kränkning|NOUN": 16.48, "trogen|ADJ": 16.47, "underteckna|VERB": 16.47, "stilla|ADV": 16.45, "invasion|NOUN": 16.43, "enhetlig|ADJ": 16.4, "not|NOUN": 16.39, "förebygga|VERB": 16.36, "lukta|VERB": 16.36, "humanitär|ADJ": 16.32, "intelligent|ADJ": 16.32, "besvär|NOUN": 16.32, "flotta|NOUN": 16.31, "turkisk|ADJ": 16.31, "mandatperiod|NOUN": 16.3, "civilisation|NOUN": 16.28, "ursäkta|VERB": 16.25, "demonstrera|VERB": 16.24, "godta|VERB": 16.24, "andas|VERB": 16.23, "böter|NOUN": 16.23, "lärdom|NOUN": 16.23, "kyla|NOUN": 16.21, "ordinarie|ADJ": 16.21, "delegation|NOUN": 16.19, "suga|VERB": 16.18, "tränare|NOUN": 16.18, "användande|NOUN": 16.17, "arbetsgrupp|NOUN": 16.17, "operatör|NOUN": 16.17, "reporter|NOUN": 16.16, "tortyr|NOUN": 16.13, "kapten|NOUN": 16.12, "forska|VERB": 16.1, "avkastning|NOUN": 16.09, "genomsnittlig|ADJ": 16.09, "jägare|NOUN": 16.09, "makthavare|NOUN": 16.06, "löjlig|ADJ": 16.04, "skönhet|NOUN": 16.04, "orimlig|ADJ": 16.03, "matematik|NOUN": 16.02, "officiellt|ADV": 16.01, "rensa|VERB": 16.0, "utvärdera|VERB": 16.0, "onekligen|ADV": 15.99, "tonåring|NOUN": 15.99, "dagsläge|NOUN": 15.98, "entreprenör|NOUN": 15.98, "kines|NOUN": 15.98, "blivande|ADJ": 15.97, "elände|NOUN": 15.96, "glida|VERB": 15.96, "stiftelse|NOUN": 15.96, "frivilligt|ADV": 15.92, "introducera|VERB": 15.92, "korrekt|ADV": 15.92, "villigt|ADV": 15.92, "friskola|NOUN": 15.89, "smula|NOUN": 15.89, "försvåra|VERB": 15.88, "kyrklig|ADJ": 15.88, "oväntad|ADJ": 15.87, "rikedom|NOUN": 15.86, "delstat|NOUN": 15.85, "gång på gång|ADV": 15.82, "illustrera|VERB": 15.82, "centralbank|NOUN": 15.81, "grannland|NOUN": 15.79, "rasist|NOUN": 15.79, "ägande|NOUN": 15.79, "förvirrad|ADJ": 15.78, "kredit|NOUN": 15.77, "rom|NOUN": 15.77, "storstad|NOUN": 15.76, "tveka|VERB": 15.76, "överföring|NOUN": 15.76, "katolik|NOUN": 15.75, "tät|ADJ": 15.75, "fotografi|NOUN": 15.74, "förare|NOUN": 15.74, "historiker|NOUN": 15.74, "misslyckande|NOUN": 15.72, "present|NOUN": 15.71, "dödsstraff|NOUN": 15.7, "evighet|NOUN": 15.68, "enighet|NOUN": 15.66, "torn|NOUN": 15.66, "stigande|ADJ": 15.66, "förkasta|VERB": 15.65, "humör|NOUN": 15.64, "hemskt|ADV": 15.63, "moment|NOUN": 15.62, "allihop (vardagl. allihopa)|PRON": 15.6, "fritid|NOUN": 15.6, "rapportering|NOUN": 15.6, "stöld|NOUN": 15.6, "konkurrenskraft|NOUN": 15.59, "psykologisk|ADJ": 15.59, "alternativt|ADV": 15.58, "direktör|NOUN": 15.58, "skeptisk|ADJ": 15.56, "bakåt|ADV": 15.54, "lapp|NOUN": 15.53, "anlita|VERB": 15.52, "avfärda|VERB": 15.52, "likadant|ADV": 15.51, "separat|ADJ": 15.5, "överensstämma|VERB": 15.49, "finansminister|NOUN": 15.48, "format|NOUN": 15.48, "ogilla|VERB": 15.48, "omvandla|VERB": 15.48, "argumentation|NOUN": 15.47, "likadan|ADJ": 15.47, "tavla|NOUN": 15.47, "kännedom|NOUN": 15.43, "programvara|NOUN": 15.43, "skattesänkning|NOUN": 15.43, "jämlikhet|NOUN": 15.42, "chefredaktör|NOUN": 15.41, "säljare|NOUN": 15.41, "duga|VERB": 15.4, "negativt|ADV": 15.4, "arkitekt|NOUN": 15.39, "livad|ADJ": 15.38, "passagerare|NOUN": 15.38, "finans|NOUN": 15.38, "ekonom|NOUN": 15.37, "läsvärd|ADJ": 15.37, "obegriplig|ADJ": 15.37, "skam|NOUN": 15.36, "skicklig|ADJ": 15.36, "störta|VERB": 15.34, "överta|VERB": 15.33, "feminist|NOUN": 15.32, "orättvisa|NOUN": 15.32, "stadsdel|NOUN": 15.32, "årligen|ADV": 15.32, "utbyggnad|NOUN": 15.32, "beskattning|NOUN": 15.29, "återge|VERB": 15.29, "koka|VERB": 15.27, "taliban|NOUN": 15.27, "skara|NOUN": 15.26, "bröllop|NOUN": 15.25, "mormor|NOUN": 15.25, "pasta|NOUN": 15.25, "itu|PART": 15.24, "fan|NOUN": 15.23, "syskon|NOUN": 15.23, "tillverkning|NOUN": 15.22, "bunden|ADJ": 15.21, "gitarr|NOUN": 15.21, "diagnos|NOUN": 15.19, "häftig|ADJ": 15.19, "överklaga|VERB": 15.19, "strejk|NOUN": 15.18, "tvång|NOUN": 15.18, "dödsfall|NOUN": 15.18, "import|NOUN": 15.18, "formellt|ADV": 15.17, "rund|ADJ": 15.17, "sambo|NOUN": 15.17, "teknologi|NOUN": 15.17, "iransk|ADJ": 15.16, "någorlunda|ADV": 15.16, "genomgång|NOUN": 15.15, "grundskola|NOUN": 15.15, "framställning|NOUN": 15.14, "rådgivare|NOUN": 15.14, "vrida|VERB": 15.14, "behaglig|ADJ": 15.13, "fästa|VERB": 15.13, "målning|NOUN": 15.13, "underskott|NOUN": 15.13, "framme|ADV": 15.11, "imperium|NOUN": 15.11, "lönsam|ADJ": 15.11, "söder|NOUN": 15.11, "successivt|ADV": 15.1, "hänvisning|NOUN": 15.1, "konsekvent|ADV": 15.1, "isolerad|ADJ": 15.09, "handlingsplan|NOUN": 15.09, "tvåa|NOUN": 15.09, "häva|VERB": 15.06, "upphäva|VERB": 15.06, "färdighet|NOUN": 15.05, "självmord|NOUN": 15.04, "svärd|NOUN": 15.04, "stall|NOUN": 15.03, "styre|NOUN": 15.01, "fristående|ADJ": 14.99, "ilska|NOUN": 14.99, "dumt|ADJ": 14.98, "offentliggöra|VERB": 14.97, "privatperson|NOUN": 14.97, "kompensera|VERB": 14.96, "överraskning|NOUN": 14.96, "stängd|ADJ": 14.94, "tröja|NOUN": 14.92, "komponent|NOUN": 14.91, "festival|NOUN": 14.9, "lågkonjunktur|NOUN": 14.89, "återställa|VERB": 14.89, "skandal|NOUN": 14.89, "med hänvisning till|ADP": 14.88, "förutse|VERB": 14.87, "minst sagt|ADV": 14.87, "stötta|VERB": 14.87, "fantastiskt|ADV": 14.85, "karl|NOUN": 14.85, "aggressiv|ADJ": 14.84, "härmed|ADV": 14.84, "avsaknad|NOUN": 14.83, "kemisk|ADJ": 14.83, "saknad|NOUN": 14.83, "raket|NOUN": 14.81, "tunnelbana|NOUN": 14.81, "värma|VERB": 14.81, "kommunistparti|NOUN": 14.79, "marginal|NOUN": 14.79, "respektive|ADV": 14.79, "gravid|ADJ": 14.78, "kniv|NOUN": 14.78, "ramla|VERB": 14.78, "villa|NOUN": 14.78, "dryg|ADJ": 14.77, "lampa|NOUN": 14.77, "överdriven|ADJ": 14.76, "back|NOUN": 14.76, "kusin|NOUN": 14.76, "knapp|NOUN": 14.75, "skynda|VERB": 14.75, "privatliv|NOUN": 14.75, "toalett|NOUN": 14.75, "bada|VERB": 14.73, "lustig|ADJ": 14.73, "provins|NOUN": 14.73, "orättvis|ADJ": 14.72, "sexualitet|NOUN": 14.72, "upptäckt|NOUN": 14.72, "kreativitet|NOUN": 14.71, "lagråd|NOUN": 14.71, "malm|NOUN": 14.68, "referera|VERB": 14.68, "teologi|NOUN": 14.68, "arkitektur|NOUN": 14.67, "förvalta|VERB": 14.67, "rättsväsende|NOUN": 14.67, "lord|NOUN": 14.66, "poet|NOUN": 14.65, "stuga|NOUN": 14.63, "regna|VERB": 14.62, "spekulera|VERB": 14.62, "bonus|NOUN": 14.6, "längtan|NOUN": 14.6, "rymd|NOUN": 14.6, "fruktansvärt|ADV": 14.58, "bad|NOUN": 14.55, "förhör|NOUN": 14.53, "likvärdig|ADJ": 14.53, "upplösa|VERB": 14.52, "blockera|VERB": 14.5, "fröken|NOUN": 14.5, "hysa|VERB": 14.49, "klipp|NOUN": 14.49, "äganderätt|NOUN": 14.49, "akademi|NOUN": 14.48, "benämna|VERB": 14.48, "indisk|ADJ": 14.48, "rosa|ADJ": 14.48, "tycke|NOUN": 14.48, "avlägsen|ADJ": 14.47, "konstigt|ADV": 14.46, "marknadsekonomi|NOUN": 14.46, "uppta|VERB": 14.46, "utland|NOUN": 14.44, "erinra|VERB": 14.43, "finanser|NOUN": 14.43, "lärande|NOUN": 14.43, "råvara|NOUN": 14.42, "förenlig|ADJ": 14.4, "klättra|VERB": 14.39, "berättigad|ADJ": 14.39, "brottsling|NOUN": 14.39, "tillhörande|ADJ": 14.37, "delaktig|ADJ": 14.36, "rusa|VERB": 14.36, "änka|NOUN": 14.35, "plugga|VERB": 14.34, "prins|NOUN": 14.34, "mystisk|ADJ": 14.33, "same|NOUN": 14.33, "bar|NOUN": 14.32, "indirekt|ADV": 14.32, "webbsida|NOUN": 14.32, "avveckla|VERB": 14.3, "bygge|NOUN": 14.3, "föredrag|NOUN": 14.3, "bibehålla|VERB": 14.29, "näring|NOUN": 14.29, "poesi|NOUN": 14.28, "smyga|VERB": 14.28, "förort|NOUN": 14.27, "genetisk|ADJ": 14.26, "sorglig|ADJ": 14.25, "fransman|NOUN": 14.25, "genre|NOUN": 14.25, "lat|ADJ": 14.25, "lastbil|NOUN": 14.23, "vårda|VERB": 14.22, "lista|VERB": 14.2, "inledande|ADJ": 14.19, "debattör|NOUN": 14.19, "premiär|NOUN": 14.18, "redskap|NOUN": 14.18, "vila|NOUN": 14.18, "novell|NOUN": 14.16, "väsentligt|ADV": 14.16, "matte|NOUN": 14.15, "anförande|NOUN": 14.12, "hyra|NOUN": 14.12, "mogen|ADJ": 14.12, "osynlig|ADJ": 14.12, "besvärlig|ADJ": 14.1, "dansk|NOUN": 14.1, "överskott|NOUN": 14.09, "kompromiss|NOUN": 14.07, "uppskattning|NOUN": 14.07, "kvart|NOUN": 14.05, "spekulation|NOUN": 14.05, "urban|ADJ": 14.05, "begriplig|ADJ": 14.04, "träff|NOUN": 14.04, "flykt|NOUN": 14.03, "poker|NOUN": 14.03, "uppgörelse|NOUN": 14.03, "besvikelse|NOUN": 14.03, "gradvis|ADV": 14.03, "acceptabel|ADJ": 14.01, "lugna|VERB": 14.01, "skräck|NOUN": 14.01, "komplett|ADJ": 14.0, "norr om|ADP": 13.99, "förhållandevis|ADV": 13.97, "hugga|VERB": 13.97, "massmedium|NOUN": 13.97, "varpå|ADV": 13.97, "åtala|VERB": 13.97, "gris|NOUN": 13.96, "medverkan|NOUN": 13.95, "märkligt|ADV": 13.95, "uppehållstillstånd|NOUN": 13.95, "original|NOUN": 13.92, "utdelning|NOUN": 13.92, "julklapp|NOUN": 13.91, "klapp|NOUN": 13.91, "långvarig|ADJ": 13.91, "still|ADV": 13.91, "sammansättning|NOUN": 13.89, "oändlig|ADJ": 13.89, "oerhörd|ADJ": 13.87, "rast|NOUN": 13.87, "skapare|NOUN": 13.87, "benämning|NOUN": 13.86, "transportera|VERB": 13.86, "uppdelning|NOUN": 13.85, "väsen|NOUN": 13.85, "islamist|NOUN": 13.84, "självklarhet|NOUN": 13.84, "beaktande|NOUN": 13.82, "i kombination med|ADP": 13.82, "reta|VERB": 13.82, "trakt|NOUN": 13.82, "inledningsvis|ADV": 13.82, "krog|NOUN": 13.82, "enig|ADJ": 13.81, "ärva|VERB": 13.81, "jätte|NOUN": 13.8, "börda|NOUN": 13.79, "föregå|VERB": 13.79, "publicering|NOUN": 13.79, "skifte|NOUN": 13.79, "aktivist|NOUN": 13.77, "guide|NOUN": 13.77, "smälta|VERB": 13.77, "styrka|VERB": 13.77, "frysa|VERB": 13.76, "noggrann|ADJ": 13.76, "systematisk|ADJ": 13.75, "tillträde|NOUN": 13.75, "oväntat|ADV": 13.72, "kompetent|ADJ": 13.7, "prostitution|NOUN": 13.7, "skick|NOUN": 13.7, "mätt|ADJ": 13.7, "inköp|NOUN": 13.68, "ficka|NOUN": 13.68, "nederlag|NOUN": 13.67, "ansökning|NOUN": 13.66, "verkligt|ADV": 13.66, "story|NOUN": 13.65, "byrå|NOUN": 13.64, "dryck|NOUN": 13.64, "smidig|ADJ": 13.64, "synvinkel|NOUN": 13.64, "så gott som|ADV": 13.64, "försvaga|VERB": 13.62, "gräs|NOUN": 13.62, "förfluten|ADJ": 13.61, "simma|VERB": 13.6, "fysik|NOUN": 13.6, "hockey|NOUN": 13.6, "produktivitet|NOUN": 13.58, "incitament|NOUN": 13.57, "kontrast|NOUN": 13.56, "läpp|NOUN": 13.56, "progressiv|ADJ": 13.56, "anmärkningsvärd|ADJ": 13.55, "mobil|NOUN": 13.55, "tull|NOUN": 13.55, "fotografera (vardagl. fota)|VERB": 13.54, "skärm|NOUN": 13.54, "databas|NOUN": 13.53, "fynd|NOUN": 13.53, "bekymmer|NOUN": 13.53, "underhåll|NOUN": 13.53, "i gång (el. igång)|ADV": 13.51, "tätt|ADV": 13.51, "överlägsen|ADJ": 13.51, "grek|NOUN": 13.5, "kedja|NOUN": 13.49, "sår|NOUN": 13.47, "uppenbarelse|NOUN": 13.47, "utfall|NOUN": 13.47, "naiv|ADJ": 13.46, "still|ADJ": 13.46, "morgondag|NOUN": 13.46, "nöd|NOUN": 13.46, "motorväg|NOUN": 13.45, "utvecklingsland|NOUN": 13.45, "avhandling|NOUN": 13.44, "godis|NOUN": 13.44, "ko|NOUN": 13.44, "påvisa|VERB": 13.44, "trampa|VERB": 13.42, "ambassadör|NOUN": 13.41, "torka|VERB": 13.41, "så att säga|ADV": 13.4, "titt|NOUN": 13.4, "spränga|VERB": 13.39, "halva|NOUN": 13.38, "känneteckna|VERB": 13.38, "ombud|NOUN": 13.38, "ortodox|ADJ": 13.37, "problematisk|ADJ": 13.37, "virus|NOUN": 13.35, "himmelsk|ADJ": 13.34, "uppsats|NOUN": 13.34, "strålande|ADJ": 13.34, "bindande|ADJ": 13.33, "alltjämt|ADV": 13.32, "jämt|ADV": 13.32, "hungrig|ADJ": 13.31, "elak|ADJ": 13.3, "bosättning|NOUN": 13.29, "miljövänlig|ADJ": 13.28, "förfogande|NOUN": 13.26, "lucka|NOUN": 13.26, "procentenhet|NOUN": 13.26, "sammanträde|NOUN": 13.26, "musikalisk|ADJ": 13.25, "självförtroende|NOUN": 13.23, "cool|ADJ": 13.21, "fördjupa|VERB": 13.21, "ingång|NOUN": 13.2, "sed|NOUN": 13.19, "taxi|NOUN": 13.19, "vänja|VERB": 13.19, "författning|NOUN": 13.18, "huvudperson|NOUN": 13.18, "hypotes|NOUN": 13.18, "panik|NOUN": 13.18, "stämma|NOUN": 13.18, "avslutning|NOUN": 13.18, "deklaration|NOUN": 13.18, "sväng|NOUN": 13.17, "presidentval|NOUN": 13.16, "undgå|VERB": 13.15, "illusion|NOUN": 13.12, "international|NOUN": 13.12, "intrång|NOUN": 13.12, "skattepengar|NOUN": 13.12, "stolthet|NOUN": 13.11, "utnyttjande|NOUN": 13.11, "överlevnad|NOUN": 13.11, "problematik|NOUN": 13.1, "sällsynt|ADJ": 13.1, "dumhet|NOUN": 13.09, "flöde|NOUN": 13.09, "jättebra|ADJ": 13.08, "i jämförelse med|ADP": 13.07, "medborgarskap|NOUN": 13.04, "snack|NOUN": 13.04, "parallellt|ADV": 13.03, "påföljd|NOUN": 13.03, "söder om|ADP": 13.02, "strax efter|ADV": 13.01, "talang|NOUN": 13.01, "varmt|ADV": 13.01, "pjäs|NOUN": 13.0, "kansli|NOUN": 12.99, "lagligt|ADV": 12.99, "sand|NOUN": 12.99, "fildelare|NOUN": 12.98, "liga|NOUN": 12.98, "parlamentarisk|ADJ": 12.98, "vittnesbörd|NOUN": 12.96, "avrätta|VERB": 12.96, "fiske|NOUN": 12.96, "gynnsam|ADJ": 12.96, "dokumentär|NOUN": 12.95, "dödlig|ADJ": 12.95, "beteckning|NOUN": 12.94, "jämte|ADP": 12.94, "uttryckligen|ADV": 12.94, "distrikt|NOUN": 12.93, "påse|NOUN": 12.93, "baksida|NOUN": 12.92, "plånbok|NOUN": 12.92, "uppsägning|NOUN": 12.92, "fullfölja|VERB": 12.91, "foga|VERB": 12.9, "psykologi|NOUN": 12.9, "hjul|NOUN": 12.89, "klänning|NOUN": 12.89, "anteckning|NOUN": 12.89, "trä|NOUN": 12.89, "belägg|NOUN": 12.88, "blunda|VERB": 12.88, "vik|NOUN": 12.88, "bråk|NOUN": 12.87, "värva|VERB": 12.87, "biblisk|ADJ": 12.86, "sikta|VERB": 12.86, "uteslutande|ADV": 12.86, "pryl|NOUN": 12.85, "begravning|NOUN": 12.84, "naturligt|ADV": 12.84, "bredd|NOUN": 12.83, "frälsning|NOUN": 12.82, "funktionshinder|NOUN": 12.82, "såvida|SCONJ": 12.82, "avvika|VERB": 12.81, "influensa|NOUN": 12.81, "medvetenhet|NOUN": 12.8, "muskel|NOUN": 12.8, "ointressant|ADJ": 12.8, "samhällelig|ADJ": 12.8, "apropå|ADP": 12.78, "cirkel|NOUN": 12.78, "rekord|NOUN": 12.78, "bemärkelse|NOUN": 12.77, "djävul|NOUN": 12.76, "tålamod|NOUN": 12.75, "utspel|NOUN": 12.75, "verkställa|VERB": 12.75, "hjälpmedel|NOUN": 12.74, "riksdagsval|NOUN": 12.74, "svära|VERB": 12.74, "tagg|NOUN": 12.74, "deklarera|VERB": 12.73, "meningsfull|ADJ": 12.73, "i anslutning till|ADP": 12.71, "rimligen|ADV": 12.71, "minut (förk. min.)|NOUN": 12.69, "annanstans|ADV": 12.68, "knapp|ADJ": 12.68, "kvartal|NOUN": 12.68, "party|NOUN": 12.68, "imponera|VERB": 12.67, "innanför|ADP": 12.67, "expansion|NOUN": 12.66, "vaken|ADJ": 12.66, "kunnig|ADJ": 12.64, "scenario|NOUN": 12.64, "leverans|NOUN": 12.62, "medelstor|ADJ": 12.62, "salt|NOUN": 12.62, "sannolik|ADJ": 12.62, "vänskap|NOUN": 12.62, "farmor|NOUN": 12.61, "tiotusentals|ADV": 12.61, "lokalt|ADV": 12.6, "frigöra|VERB": 12.59, "prestation|NOUN": 12.59, "olämplig|ADJ": 12.58, "belöning|NOUN": 12.57, "styrning|NOUN": 12.57, "säte|NOUN": 12.57, "sjukförsäkring|NOUN": 12.56, "upplysa|VERB": 12.56, "halvtimme|NOUN": 12.55, "uppsättning|NOUN": 12.54, "sms|NOUN": 12.54, "elektrisk|ADJ": 12.53, "folkbildning|NOUN": 12.53, "kriminalitet|NOUN": 12.53, "födelse|NOUN": 12.52, "registrering|NOUN": 12.52, "nord|NOUN": 12.5, "färdas|VERB": 12.5, "världsbild|NOUN": 12.49, "brista|VERB": 12.48, "prinsessa|NOUN": 12.48, "överlåta|VERB": 12.48, "konsumera|VERB": 12.47, "vardaglig|ADJ": 12.47, "besättning|NOUN": 12.46, "manus|NOUN": 12.46, "mestadels|ADV": 12.46, "glädjande|ADJ": 12.46, "imperialism|NOUN": 12.46, "departement|NOUN": 12.44, "förfölja|VERB": 12.44, "operativ|ADJ": 12.44, "fullmäktige|NOUN": 12.42, "kommunfullmäktige|NOUN": 12.42, "nyliberal|ADJ": 12.39, "sparande|NOUN": 12.39, "interpellation|NOUN": 12.39, "marxism|NOUN": 12.39, "trång|ADJ": 12.39, "angelägenhet|NOUN": 12.38, "potatis|NOUN": 12.38, "medeltida|ADJ": 12.37, "underhållande|ADJ": 12.37, "ensamhet|NOUN": 12.36, "noggrant|ADV": 12.36, "sprit|NOUN": 12.36, "panna|NOUN": 12.35, "sakfråga|NOUN": 12.34, "brun|ADJ": 12.33, "kind|NOUN": 12.33, "förekomst|NOUN": 12.32, "härifrån|ADV": 12.32, "okunnig|ADJ": 12.32, "oförändrad|ADJ": 12.32, "sedermera|ADV": 12.31, "möjligtvis|ADV": 12.3, "fordra|VERB": 12.29, "förhållningssätt|NOUN": 12.29, "hall|NOUN": 12.29, "regelbunden|ADJ": 12.28, "klassiker|NOUN": 12.27, "uppkomst|NOUN": 12.27, "vägledning|NOUN": 12.27, "kika|VERB": 12.26, "dos|NOUN": 12.25, "försiktigt|ADV": 12.25, "blodig|ADJ": 12.25, "dynamisk|ADJ": 12.25, "portion|NOUN": 12.25, "smutsig|ADJ": 12.25, "svika|VERB": 12.24, "smått|ADV": 12.23, "bortsett från|ADP": 12.22, "förstärkning|NOUN": 12.22, "förteckning|NOUN": 12.22, "narkotikum|NOUN": 12.21, "björn|NOUN": 12.2, "engelsman|NOUN": 12.2, "utropa|VERB": 12.2, "fascism|NOUN": 12.19, "gnälla|VERB": 12.19, "underbart|ADV": 12.19, "ankomst|NOUN": 12.18, "barnbarn|NOUN": 12.18, "gudstjänst|NOUN": 12.18, "pott|NOUN": 12.18, "regissör|NOUN": 12.18, "turk|NOUN": 12.18, "hylla|NOUN": 12.18, "tillfälligt|ADV": 12.18, "ungdomsförbund|NOUN": 12.16, "eftersträva|VERB": 12.15, "förflytta|VERB": 12.15, "sekreterare|NOUN": 12.15, "missnöjd|ADJ": 12.14, "värdelös|ADJ": 12.13, "doft|NOUN": 12.12, "passiv|ADJ": 12.11, "uppfinning|NOUN": 12.11, "språklig|ADJ": 12.1, "härska|VERB": 12.1, "kast|NOUN": 12.1, "sympati|NOUN": 12.1, "behörighet|NOUN": 12.09, "förknippa|VERB": 12.09, "insändare|NOUN": 12.09, "judendom|NOUN": 12.09, "sjuksköterska|NOUN": 12.07, "tält|NOUN": 12.07, "uppgång|NOUN": 12.07, "inskränka|VERB": 12.06, "prestera|VERB": 12.06, "udda|ADJ": 12.06, "journal|NOUN": 12.06, "diplomatisk|ADJ": 12.05, "tillfredsställande|ADJ": 12.04, "förakt|NOUN": 12.03, "regera|VERB": 12.03, "indirekt|ADJ": 12.01, "gyllene|ADJ": 12.0, "söderut|ADV": 12.0, "kapitalist|NOUN": 11.99, "genomslag|NOUN": 11.98, "teologisk|ADJ": 11.98, "matta|NOUN": 11.96, "medelklass|NOUN": 11.95, "målgrupp|NOUN": 11.95, "sortera|VERB": 11.95, "säkerhetspolitik|NOUN": 11.95, "födelsedag|NOUN": 11.94, "misshandla|VERB": 11.94, "mynt|NOUN": 11.94, "rörlig|ADJ": 11.94, "gods|NOUN": 11.93, "beredning|NOUN": 11.92, "traditionellt|ADV": 11.92, "bliva|VERB": 11.91, "agent|NOUN": 11.9, "exklusiv|ADJ": 11.9, "handlande|NOUN": 11.9, "socker|NOUN": 11.9, "upplopp|NOUN": 11.9, "kaka|NOUN": 11.89, "kollektivtrafik|NOUN": 11.89, "anlägga|VERB": 11.89, "upphandling|NOUN": 11.89, "breda|VERB": 11.88, "realitet|NOUN": 11.88, "marknadsföra|VERB": 11.87, "vitt|ADV": 11.87, "vrede|NOUN": 11.87, "satan|NOUN": 11.87, "statistisk|ADJ": 11.86, "ödmjuk|ADJ": 11.86, "i natt|ADV": 11.85, "klarhet|NOUN": 11.85, "långsiktigt|ADV": 11.85, "anstränga|VERB": 11.83, "generös|ADJ": 11.82, "mellanrum|NOUN": 11.82, "sken|NOUN": 11.82, "upplösning|NOUN": 11.82, "vistelse|NOUN": 11.82, "växla|VERB": 11.82, "strukturell|ADJ": 11.81, "förvärva|VERB": 11.78, "regi|NOUN": 11.78, "anka|NOUN": 11.78, "redogörelse|NOUN": 11.77, "statsmakt|NOUN": 11.77, "etta|NOUN": 11.76, "relativ|ADJ": 11.76, "vindkraft|NOUN": 11.76, "imperialistisk|ADJ": 11.75, "måltid|NOUN": 11.75, "till synes|ADV": 11.75, "belöna|VERB": 11.74, "importera|VERB": 11.74, "liter|NOUN": 11.74, "rentav|ADV": 11.74, "stormakt|NOUN": 11.74, "samtida|ADJ": 11.73, "legal|ADJ": 11.72, "principiell|ADJ": 11.72, "valfrihet|NOUN": 11.72, "tydlighet|NOUN": 11.71, "växthusgas|NOUN": 11.71, "evenemang|NOUN": 11.69, "lösenord|NOUN": 11.68, "dialekt|NOUN": 11.67, "behärska|VERB": 11.66, "föregångare|NOUN": 11.66, "homosexualitet|NOUN": 11.66, "seg|ADJ": 11.66, "licens|NOUN": 11.65, "platt|ADJ": 11.65, "iver|NOUN": 11.64, "resenär|NOUN": 11.63, "utrota|VERB": 11.63, "uppfinna|VERB": 11.62, "cup|NOUN": 11.61, "omvänd|ADJ": 11.61, "dagordning|NOUN": 11.61, "perfekt|ADV": 11.6, "splittring|NOUN": 11.6, "inbilla|VERB": 11.59, "avge|VERB": 11.58, "partnerskap|NOUN": 11.58, "löna sig|VERB": 11.57, "brutal|ADJ": 11.56, "konstruera|VERB": 11.56, "ärlighet|NOUN": 11.56, "bekväm|ADJ": 11.54, "presskonferens|NOUN": 11.54, "osannolik|ADJ": 11.53, "totalitär|ADJ": 11.53, "åtgärda|VERB": 11.53, "flickvän|NOUN": 11.53, "norrut|ADV": 11.53, "arbetstillfälle|NOUN": 11.52, "inträde|NOUN": 11.52, "släpa|VERB": 11.52, "övervägande|NOUN": 11.52, "skilsmässa|NOUN": 11.51, "utforska|VERB": 11.5, "bildande|ADJ": 11.47, "tyngd|NOUN": 11.47, "frälsare|NOUN": 11.46, "invadera|VERB": 11.46, "personuppgift|NOUN": 11.46, "förhand|NOUN": 11.46, "gruppering|NOUN": 11.46, "tekniskt|ADV": 11.46, "dagstidning|NOUN": 11.45, "oacceptabel|ADJ": 11.45, "serb|NOUN": 11.45, "flytande|ADJ": 11.45, "justera|VERB": 11.44, "adel|NOUN": 11.43, "konsult|NOUN": 11.43, "nervös|ADJ": 11.43, "sekt|NOUN": 11.42, "slöja|NOUN": 11.42, "välkommen|INTJ": 11.42, "läcka|VERB": 11.41, "afton|NOUN": 11.4, "introduktion|NOUN": 11.4, "livstid|NOUN": 11.4, "demonstrant|NOUN": 11.39, "flexibilitet|NOUN": 11.39, "hed|NOUN": 11.39, "kol|NOUN": 11.39, "uppväxt|NOUN": 11.39, "efterlysa|VERB": 11.37, "grönsak|NOUN": 11.37, "samordna|VERB": 11.37, "järn|NOUN": 11.35, "distribution|NOUN": 11.34, "automatisk|ADJ": 11.32, "transaktion|NOUN": 11.32, "däck|NOUN": 11.31, "observation|NOUN": 11.31, "typiskt|ADV": 11.31, "inskränkning|NOUN": 11.3, "mata|VERB": 11.3, "paradis|NOUN": 11.3, "ingenjör|NOUN": 11.29, "koncentration|NOUN": 11.29, "plus|NOUN": 11.29, "dugg|NOUN": 11.27, "samtid|NOUN": 11.27, "uppståndelse|NOUN": 11.27, "slaveri|NOUN": 11.26, "ålägga|VERB": 11.26, "framkalla|VERB": 11.25, "utkast|NOUN": 11.25, "framträdande|ADJ": 11.25, "desperat|ADJ": 11.25, "någon som helst|DET": 11.25, "flitigt|ADV": 11.22, "offensiv|NOUN": 11.22, "sångare|NOUN": 11.22, "ingrepp|NOUN": 11.21, "otalig|ADJ": 11.21, "diagram|NOUN": 11.2, "inbjuda|VERB": 11.2, "motivation|NOUN": 11.2, "utplåna|VERB": 11.2, "gymnasieskola|NOUN": 11.19, "bearbeta|VERB": 11.18, "förlåtelse|NOUN": 11.18, "snurra|VERB": 11.18, "skildring|NOUN": 11.18, "sändning|NOUN": 11.18, "baby|NOUN": 11.18, "förvara|VERB": 11.17, "rabatt|NOUN": 11.17, "rota|VERB": 11.17, "apa|NOUN": 11.16, "sammanställa|VERB": 11.16, "stirra|VERB": 11.16, "avgörande|NOUN": 11.15, "manifestation|NOUN": 11.15, "uppenbara|VERB": 11.15, "maila|VERB": 11.14, "medmänniska|NOUN": 11.14, "genombrott|NOUN": 11.12, "proletär|ADJ": 11.12, "fika|NOUN": 11.1, "spaning|NOUN": 11.1, "beordra|VERB": 11.1, "förbinda|VERB": 11.1, "jämförbar|ADJ": 11.1, "socialt|ADV": 11.1, "fullgöra|VERB": 11.09, "förr eller senare|ADV": 11.09, "palm|NOUN": 11.08, "förvirring|NOUN": 11.08, "privatisering|NOUN": 11.08, "chock|NOUN": 11.07, "oundviklig|ADJ": 11.06, "samtycke|NOUN": 11.06, "förband|NOUN": 11.04, "missbruka|VERB": 11.03, "förvärra|VERB": 11.02, "investerare|NOUN": 11.02, "vackert|ADV": 11.02, "utbredd|ADJ": 11.02, "bio|NOUN": 11.01, "oförmåga|NOUN": 11.01, "sammanlagd|ADJ": 11.0, "klippa|NOUN": 11.0, "cd|NOUN": 10.99, "knut|NOUN": 10.98, "fras|NOUN": 10.97, "indikera|VERB": 10.97, "vardera|PRON": 10.97, "arrangör|NOUN": 10.96, "profetia|NOUN": 10.96, "därutöver|ADV": 10.96, "förnya|VERB": 10.96, "hederlig|ADJ": 10.95, "inhämta|VERB": 10.95, "skånsk|ADJ": 10.95, "abstrakt|ADJ": 10.94, "dämpa|VERB": 10.94, "tillhörighet|NOUN": 10.94, "möbel|NOUN": 10.93, "ringa|ADJ": 10.93, "sky|NOUN": 10.93, "anvisning|NOUN": 10.91, "hatt|NOUN": 10.9, "tokig|ADJ": 10.9, "förvärv|NOUN": 10.89, "med flera (förk. m.fl., m fl)|ADV": 10.89, "omgående|ADV": 10.89, "bedrägeri|NOUN": 10.89, "mobilisera|VERB": 10.89, "signatur|NOUN": 10.88, "skälig|ADJ": 10.88, "expandera|VERB": 10.87, "förkunna|VERB": 10.87, "böja|VERB": 10.86, "förenkla|VERB": 10.86, "viga|VERB": 10.85, "justitieminister|NOUN": 10.84, "fjärdedel|NOUN": 10.83, "substans|NOUN": 10.83, "tömma|VERB": 10.83, "utmärka|VERB": 10.83, "ende|ADJ": 10.82, "förnyelse|NOUN": 10.82, "subjektiv|ADJ": 10.82, "burk|NOUN": 10.81, "human|ADJ": 10.81, "mista|VERB": 10.81, "sanktion|NOUN": 10.81, "fler och fler|PRON": 10.8, "omsättning|NOUN": 10.8, "besitta|VERB": 10.78, "initiera|VERB": 10.78, "skrivande|NOUN": 10.77, "hänseende|NOUN": 10.76, "härstamma|VERB": 10.76, "censur|NOUN": 10.75, "kollektiv|NOUN": 10.75, "promenera|VERB": 10.75, "supa|VERB": 10.75, "legitimitet|NOUN": 10.75, "befäl|NOUN": 10.74, "sökande|NOUN": 10.65, "pojkvän|NOUN": 10.71, "poängtera|VERB": 10.71, "överträdelse|NOUN": 10.71, "klimatfråga|NOUN": 10.7, "telefonsamtal|NOUN": 10.7, "beredskap|NOUN": 10.68, "vers|NOUN": 10.68, "monarki|NOUN": 10.67, "ockupera|VERB": 10.67, "skum|ADJ": 10.67, "turism|NOUN": 10.67, "befrielse|NOUN": 10.65, "byxa|NOUN": 10.65, "rekrytera|VERB": 10.65, "förmögenhet|NOUN": 10.64, "gången|ADJ": 10.64, "liksom|SCONJ": 10.64, "äpple|NOUN": 10.64, "höjdpunkt|NOUN": 10.63, "sammanställning|NOUN": 10.62, "underhållning|NOUN": 10.62, "uppbyggnad|NOUN": 10.62, "etablissemang|NOUN": 10.61, "kontinuerligt|ADV": 10.61, "krama|VERB": 10.61, "missförstånd|NOUN": 10.61, "nationalistisk|ADJ": 10.61, "obalans|NOUN": 10.61, "nyår|NOUN": 10.61, "produktiv|ADJ": 10.6, "till rätta|ADV": 10.6, "avveckling|NOUN": 10.59, "provocera|VERB": 10.59, "erfaren|ADJ": 10.58, "blank|ADJ": 10.58, "singel|NOUN": 10.58, "försörjning|NOUN": 10.55, "irländsk|ADJ": 10.55, "kurd|NOUN": 10.55, "psykolog|NOUN": 10.55, "samtala|VERB": 10.55, "sekel|NOUN": 10.55, "federal|ADJ": 10.54, "frustration|NOUN": 10.54, "fundamental|ADJ": 10.54, "omge|VERB": 10.54, "företa|VERB": 10.53, "utdrag|NOUN": 10.53, "fram och tillbaka|ADV": 10.53, "lågt|ADV": 10.53, "skal|NOUN": 10.53, "irakisk|ADJ": 10.52, "parallell|NOUN": 10.52, "avslag|NOUN": 10.51, "emellanåt|ADV": 10.51, "källare|NOUN": 10.51, "merpart|NOUN": 10.51, "vetskap|NOUN": 10.51, "delägare|NOUN": 10.5, "distans|NOUN": 10.5, "eliminera|VERB": 10.5, "i motsats till|ADP": 10.5, "tolerans|NOUN": 10.5, "krigare|NOUN": 10.49, "bosätta|VERB": 10.49, "filma|VERB": 10.48, "upplägg|NOUN": 10.48, "föda|NOUN": 10.47, "överläggning|NOUN": 10.47, "miss|NOUN": 10.46, "moské|NOUN": 10.46, "passion|NOUN": 10.46, "zon|NOUN": 10.46, "tunga|NOUN": 10.45, "vass|ADJ": 10.45, "klient|NOUN": 10.44, "spana|VERB": 10.44, "utbetalning|NOUN": 10.44, "obetydlig|ADJ": 10.43, "kurdisk|ADJ": 10.42, "relevans|NOUN": 10.41, "förutsatt att|SCONJ": 10.4, "motarbeta|VERB": 10.4, "påtryckning|NOUN": 10.4, "efterföljande|ADJ": 10.39, "nyhetsbrev|NOUN": 10.39, "årsskifte|NOUN": 10.39, "avvikelse|NOUN": 10.39, "tilltala|VERB": 10.39, "stift|NOUN": 10.38, "hemlös|ADJ": 10.37, "splittra|VERB": 10.37, "bosätta sig|VERB": 10.36, "bekräftelse|NOUN": 10.35, "försvarsminister|NOUN": 10.35, "dokumentera|VERB": 10.34, "lydnad|NOUN": 10.34, "tragedi|NOUN": 10.34, "organism|NOUN": 10.33, "socialtjänst|NOUN": 10.33, "tillskriva|VERB": 10.33, "humanist|NOUN": 10.32, "snett|ADV": 10.32, "firma|NOUN": 10.32, "förankring|NOUN": 10.32, "reporänta|NOUN": 10.32, "sekulär|ADJ": 10.31, "fortsättningsvis|ADV": 10.3, "erfara|VERB": 10.29, "inblandning|NOUN": 10.29, "signalspaning|NOUN": 10.29, "svininfluensa|NOUN": 10.29, "liknelse|NOUN": 10.28, "beväpnad|ADJ": 10.28, "härligt|ADV": 10.27, "ingripande|NOUN": 10.26, "pigg|ADJ": 10.25, "bebyggelse|NOUN": 10.25, "fysiskt|ADV": 10.25, "romantisk|ADJ": 10.25, "ingående|ADJ": 10.24, "märkning|NOUN": 10.24, "lojalitet|NOUN": 10.23, "penna|NOUN": 10.23, "får|NOUN": 10.22, "illustration|NOUN": 10.22, "rock|NOUN": 10.22, "innehav|NOUN": 10.21, "tilltro|NOUN": 10.2, "dvd|NOUN": 10.18, "bensin|NOUN": 10.18, "bromsa|VERB": 10.18, "bråka|VERB": 10.18, "kula|NOUN": 10.18, "svält|NOUN": 10.18, "klo|NOUN": 10.18, "sektion|NOUN": 10.18, "avskaffande|NOUN": 10.17, "examen|NOUN": 10.17, "religionsfrihet|NOUN": 10.16, "utåt|ADV": 10.16, "balansera|VERB": 10.15, "heltid|NOUN": 10.15, "hemifrån|ADV": 10.15, "stifta|VERB": 10.15, "verkställande|ADJ": 10.15, "asyl|NOUN": 10.13, "graviditet|NOUN": 10.13, "korsa|VERB": 10.13, "avlägsna|VERB": 10.12, "beställning|NOUN": 10.12, "fasad|NOUN": 10.12, "infinna sig|VERB": 10.12, "hyfsat|ADV": 10.11, "julafton|NOUN": 10.11, "organisk|ADJ": 10.11, "åtnjuta|VERB": 10.11, "för alltid|ADV": 10.11, "hemmaplan|NOUN": 10.1, "kloster|NOUN": 10.1, "förlita sig|VERB": 10.09, "förlägga|VERB": 10.09, "spontan|ADJ": 10.09, "informell|ADJ": 10.08, "förvåning|NOUN": 10.07, "iaktta|VERB": 10.07, "körkort|NOUN": 10.07, "försäkringsbolag|NOUN": 10.06, "missnöje|NOUN": 10.05, "etnicitet|NOUN": 10.04, "inbjudan|NOUN": 10.03, "dyster|ADJ": 10.03, "okunskap|NOUN": 10.03, "garanterat|ADV": 10.02, "sammanfattningsvis|ADV": 10.02, "spark|NOUN": 10.02, "arbetsdag|NOUN": 10.01, "silver|NOUN": 10.01, "organisatorisk|ADJ": 10.0, "slutgiltig|ADJ": 10.0, "tungt|ADV": 10.0, "bekänna|VERB": 9.99, "kostym|NOUN": 9.99, "schema|NOUN": 9.99, "långtgående|ADJ": 9.98, "mask|NOUN": 9.98, "materiel|NOUN": 9.98, "mobbning|NOUN": 9.98, "leksak|NOUN": 9.96, "spridd|ADJ": 9.96, "stava|VERB": 9.96, "tillit|NOUN": 9.96, "modig|ADJ": 9.95, "utbrott|NOUN": 9.95, "apparat|NOUN": 9.94, "disk|NOUN": 9.92, "drama|NOUN": 9.92, "exportera|VERB": 9.92, "försoning|NOUN": 9.92, "universell|ADJ": 9.92, "beroende|NOUN": 9.91, "surfa|VERB": 9.91, "diktator|NOUN": 9.9, "passage|NOUN": 9.9, "inbyggd|ADJ": 9.9, "plåga|VERB": 9.89, "strikt|ADJ": 9.88, "utlova|VERB": 9.88, "riksbank|NOUN": 9.87, "återta|VERB": 9.87, "dokumentation|NOUN": 9.86, "ingrediens|NOUN": 9.86, "inträda|VERB": 9.86, "show|NOUN": 9.86, "bak|ADV": 9.84, "delaktighet|NOUN": 9.84, "i viss mån|ADV": 9.83, "odling|NOUN": 9.83, "vardagsrum|NOUN": 9.83, "fascinerande|ADJ": 9.82, "kontext|NOUN": 9.82, "lina|NOUN": 9.81, "folkhögskola|NOUN": 9.79, "glasögon|NOUN": 9.79, "inviga|VERB": 9.79, "rop|NOUN": 9.79, "varannan|DET": 9.79, "disciplin|NOUN": 9.77, "europé|NOUN": 9.77, "härskare|NOUN": 9.77, "återkomst|NOUN": 9.77, "i fred|ADV": 9.76, "kompensation|NOUN": 9.75, "representativ|ADJ": 9.75, "strömma|VERB": 9.75, "kartlägga|VERB": 9.75, "systematiskt|ADV": 9.74, "i relation till|ADP": 9.73, "uppe|PART": 9.73, "yxa|NOUN": 9.73, "bevakning|NOUN": 9.72, "missionär|NOUN": 9.72, "rätta|NOUN": 9.72, "bekännelse|NOUN": 9.71, "ensidig|ADJ": 9.71, "högtid|NOUN": 9.71, "institutionell|ADJ": 9.71, "psykiskt|ADV": 9.71, "skjorta|NOUN": 9.71, "under förutsättning att|SCONJ": 9.71, "rehabilitering|NOUN": 9.7, "skärgård|NOUN": 9.7, "övervinna|VERB": 9.7, "enkät|NOUN": 9.69, "garderob|NOUN": 9.69, "läxa|NOUN": 9.69, "med avseende på|ADP": 9.69, "trumma|NOUN": 9.68, "pol|NOUN": 9.68, "choklad|NOUN": 9.67, "återhämtning|NOUN": 9.67, "bakterie|NOUN": 9.65, "exploatering|NOUN": 9.65, "kärnkraftverk|NOUN": 9.65, "stig|NOUN": 9.65, "primär|ADJ": 9.64, "republikan|NOUN": 9.64, "gestalt|NOUN": 9.63, "konstitutionell|ADJ": 9.63, "avslutningsvis|ADV": 9.62, "indian|NOUN": 9.62, "ingenstans|ADV": 9.61, "nuförtiden (el. nu för tiden)|ADV": 9.61, "runda|NOUN": 9.6, "baltisk|ADJ": 9.59, "farfar|NOUN": 9.59, "förtydliga|VERB": 9.59, "gärningsman|NOUN": 9.59, "succé|NOUN": 9.59, "tröst|NOUN": 9.59, "epok|NOUN": 9.58, "intention|NOUN": 9.58, "nedskärning|NOUN": 9.58, "tillika|ADV": 9.58, "remiss|NOUN": 9.57, "skåda|VERB": 9.57, "bevittna|VERB": 9.56, "främling|NOUN": 9.56, "juridik|NOUN": 9.56, "utvisning|NOUN": 9.56, "folkrätt|NOUN": 9.55, "legitim|ADJ": 9.55, "bostadsområde|NOUN": 9.54, "egyptisk|ADJ": 9.54, "glatt|ADV": 9.54, "hyresgäst|NOUN": 9.54, "radikalt|ADV": 9.54, "vinge|NOUN": 9.54, "klassa|VERB": 9.53, "legend|NOUN": 9.53, "öre|NOUN": 9.52, "nazistisk|ADJ": 9.51, "varsin|PRON": 9.51, "begrava|VERB": 9.5, "funktionsnedsättning|NOUN": 9.5, "kontra|ADP": 9.5, "persisk|ADJ": 9.49, "tillskott|NOUN": 9.48, "klagomål|NOUN": 9.47, "konstverk|NOUN": 9.47, "kortsiktig|ADJ": 9.47, "avliden|ADJ": 3.27, "backe|NOUN": 9.46, "förespråkare|NOUN": 9.46, "indikator|NOUN": 9.46, "nutida|ADJ": 9.46, "textstorlek|NOUN": 9.46, "åta|VERB": 9.46, "asiatisk|ADJ": 9.45, "meny|NOUN": 9.45, "muntlig|ADJ": 9.45, "nedre|ADJ": 9.45, "regeringsform|NOUN": 9.45, "otrevlig|ADJ": 9.44, "publikation|NOUN": 9.44, "halt|NOUN": 9.43, "borg|NOUN": 9.42, "pedofil|NOUN": 9.42, "porträtt|NOUN": 9.42, "utomstående|ADJ": 9.42, "ironi|NOUN": 9.4, "manipulera|VERB": 9.4, "afghansk|ADJ": 9.39, "jag|NOUN": 9.39, "utomhus|ADV": 9.39, "privilegium|NOUN": 9.39, "rensning|NOUN": 9.38, "etapp|NOUN": 9.37, "minimera|VERB": 9.36, "till fullo|ADV": 9.36, "representation|NOUN": 9.35, "latin|NOUN": 9.34, "måhända|ADV": 9.32, "serbisk|ADJ": 9.32, "estetisk|ADJ": 9.31, "explodera|VERB": 9.31, "folkrörelse|NOUN": 9.31, "grundare|NOUN": 9.31, "konspiration|NOUN": 9.31, "kritiskt|ADV": 9.31, "kurva|NOUN": 9.31, "operera|VERB": 9.3, "turné|NOUN": 9.3, "åskådare|NOUN": 9.29, "forntid|NOUN": 9.29, "alliansregering|NOUN": 9.28, "framgångsrikt|ADV": 9.28, "ovan|ADP": 9.28, "robot|NOUN": 9.28, "försvarare|NOUN": 9.27, "landslag|NOUN": 9.27, "proportion|NOUN": 9.27, "verkstad|NOUN": 9.27, "ask|NOUN": 9.26, "bomba|VERB": 9.26, "jeans|NOUN": 9.26, "jordbävning|NOUN": 9.26, "ratt|NOUN": 9.25, "brant|ADJ": 9.25, "befälhavare|NOUN": 9.25, "bot|NOUN": 9.25, "dusch|NOUN": 9.25, "konsensus|NOUN": 9.25, "könsneutral|ADJ": 9.25, "våldta|VERB": 9.24, "skruva|VERB": 9.22, "slutföra|VERB": 9.21, "återspegla|VERB": 9.21, "eko|NOUN": 9.2, "horisont|NOUN": 9.2, "inkomma|VERB": 9.19, "ministerråd|NOUN": 9.19, "beslutsfattare|NOUN": 9.18, "suck|NOUN": 9.18, "utlösa|VERB": 9.18, "flygbolag|NOUN": 9.18, "spegel|NOUN": 9.18, "konventionell|ADJ": 9.17, "metall|NOUN": 9.17, "återstående|ADJ": 9.17, "i fjol|ADV": 9.16, "lönsamhet|NOUN": 9.16, "vari|ADV": 9.16, "balanserad|ADJ": 9.15, "antiken|NOUN": 9.15, "innovativ|ADJ": 9.15, "utnämna|VERB": 9.15, "islamistisk|ADJ": 9.14, "pricka|VERB": 9.14, "tunnel|NOUN": 9.13, "avreglering|NOUN": 9.12, "bristfällig|ADJ": 9.12, "ensamstående|ADJ": 9.12, "inomhus|ADV": 9.12, "kapabel|ADJ": 9.12, "autonom|ADJ": 9.11, "mekanisk|ADJ": 9.11, "övertygande|ADJ": 9.11, "kvarvarande|ADJ": 9.1, "vägnar|NOUN": 9.1, "befara|VERB": 9.09, "beundra|VERB": 9.09, "förfall|NOUN": 9.09, "toppmöte|NOUN": 9.08, "trakasseri|NOUN": 9.08, "kupp|NOUN": 9.07, "bistå|VERB": 9.06, "sno|VERB": 9.06, "genuin|ADJ": 9.05, "nuläge|NOUN": 9.05, "ros|NOUN": 9.05, "tittare|NOUN": 9.05, "trasig|ADJ": 9.05, "check|NOUN": 9.04, "irrelevant|ADJ": 9.04, "moraliskt|ADV": 9.04, "överlag|ADV": 9.04, "förstånd|NOUN": 9.03, "blockad|NOUN": 9.03, "nutid|NOUN": 9.03, "omställning|NOUN": 9.03, "rumpa|NOUN": 9.02, "förebyggande|ADJ": 9.01, "notis|NOUN": 9.01, "mejl|NOUN": 9.0, "moms|NOUN": 9.0, "samspel|NOUN": 9.0, "aktiebolag|NOUN": 8.99, "jävel|NOUN": 8.99, "ledighet|NOUN": 8.99, "prat|NOUN": 8.99, "uppför|ADP": 8.99, "riksdagsbeslut|NOUN": 8.98, "balkong|NOUN": 8.97, "glass|NOUN": 8.97, "kallelse|NOUN": 8.97, "omsätta|VERB": 8.97, "destruktiv|ADJ": 8.96, "för|NOUN": 8.96, "sy|VERB": 8.96, "virtuell|ADJ": 8.96, "ärkebiskop|NOUN": 8.96, "invända|VERB": 8.95, "restriktion|NOUN": 8.95, "snar|ADJ": 8.95, "upprörd|ADJ": 8.95, "koncern|NOUN": 8.94, "minimal|ADJ": 8.94, "konvent|NOUN": 8.93, "fientlig|ADJ": 8.93, "förfader|NOUN": 8.93, "underhålla|VERB": 8.93, "vansinnig|ADJ": 8.93, "biografi|NOUN": 8.92, "räddning|NOUN": 8.92, "rör|NOUN": 8.92, "fiska|VERB": 8.91, "försämring|NOUN": 8.9, "mode|NOUN": 8.89, "programledare|NOUN": 8.89, "ytlig|ADJ": 8.89, "genomgående|ADJ": 8.88, "tron|NOUN": 8.88, "efternamn|NOUN": 8.87, "hämnd|NOUN": 8.86, "puls|NOUN": 8.86, "tidsperiod|NOUN": 8.85, "medelålder|NOUN": 8.84, "nyfikenhet|NOUN": 8.84, "barnomsorg|NOUN": 8.83, "ggr (gånger)|NOUN": 8.83, "framstående|ADJ": 8.82, "innehavare|NOUN": 8.82, "funktionshindrad|ADJ": 8.82, "isolering|NOUN": 8.82, "kreditkort|NOUN": 8.82, "otillräcklig|ADJ": 8.82, "arbetsmiljö|NOUN": 8.81, "fusk|NOUN": 8.81, "lik|NOUN": 8.81, "nationalitet|NOUN": 8.81, "smör|NOUN": 8.81, "tillträda|VERB": 8.81, "bänk|NOUN": 8.8, "korthet|NOUN": 8.8, "kungarike|NOUN": 8.8, "målvakt|NOUN": 8.8, "svans|NOUN": 8.8, "utvisa|VERB": 8.8, "lite grann|ADV": 8.79, "efterträdare|NOUN": 8.78, "närstående|ADJ": 8.78, "parallell|ADJ": 8.78, "plötslig|ADJ": 8.78, "rök|NOUN": 8.78, "skälla|VERB": 8.78, "valp|NOUN": 8.78, "fruktan|NOUN": 8.76, "rekrytering|NOUN": 8.76, "förövare|NOUN": 8.75, "popularitet|NOUN": 8.75, "symbolisera|VERB": 8.75, "kollaps|NOUN": 8.75, "kändis|NOUN": 8.74, "ont|NOUN": 8.74, "termin|NOUN": 8.74, "tills vidare|ADV": 8.74, "dilemma|NOUN": 8.73, "smärtsam|ADJ": 8.73, "holländsk|ADJ": 8.72, "klämma|VERB": 8.71, "ateist|NOUN": 8.7, "fotnot|NOUN": 8.7, "samverka|VERB": 8.7, "antik|ADJ": 8.69, "krånglig|ADJ": 8.69, "förpackning|NOUN": 8.68, "överskrida|VERB": 8.68, "aktivera|VERB": 8.68, "flytt|NOUN": 8.68, "vida|ADV": 8.68, "älg|NOUN": 8.68, "förstörelse|NOUN": 8.67, "elegant|ADJ": 8.66, "avgång|NOUN": 8.66, "montera|VERB": 8.65, "polisman|NOUN": 8.65, "preliminär|ADJ": 8.65, "primitiv|ADJ": 8.65, "avrättning|NOUN": 8.64, "nedåt|ADV": 8.64, "real|ADJ": 8.64, "överväldigande|ADJ": 8.64, "gym|NOUN": 8.63, "federation|NOUN": 8.62, "mötesplats|NOUN": 8.62, "öster|NOUN": 8.62, "beslutsfattande|NOUN": 8.61, "psykiatri|NOUN": 8.61, "handläggning|NOUN": 8.61, "utbryta|VERB": 8.61, "fientlighet|NOUN": 8.6, "inredning|NOUN": 8.6, "troll|NOUN": 8.6, "identisk|ADJ": 8.59, "riksförbund|NOUN": 8.59, "sal|NOUN": 8.59, "förtjust|ADV": 8.58, "generalsekreterare|NOUN": 8.58, "genomsyra|VERB": 8.58, "öppning|NOUN": 8.58, "obefintlig|ADJ": 8.57, "tillförlitlig|ADJ": 8.57, "näringsminister|NOUN": 8.55, "protein|NOUN": 8.55, "applåd|NOUN": 8.54, "ersättare|NOUN": 8.54, "onödigt|ADV": 8.54, "tjänstgöra|VERB": 8.54, "fastslå|VERB": 8.53, "slut|ADJ": 8.53, "solig|ADJ": 8.53, "gåta|NOUN": 8.53, "härlighet|NOUN": 8.53, "återuppta|VERB": 8.53, "fördriva|VERB": 8.52, "hertig|NOUN": 8.52, "påsk|NOUN": 8.52, "komplement|NOUN": 8.51, "modersmål|NOUN": 8.51, "beröm|NOUN": 8.5, "frö|NOUN": 8.5, "installation|NOUN": 8.5, "släcka|VERB": 8.49, "odds|NOUN": 8.48, "årsmöte|NOUN": 8.48, "arm|ADJ": 8.47, "kommunstyrelse|NOUN": 8.47, "mångkulturell|ADJ": 8.47, "varaktig|ADJ": 8.47, "horn|NOUN": 8.47, "sedel|NOUN": 8.46, "valsedel|NOUN": 8.46, "merit|NOUN": 8.46, "skinn|NOUN": 8.45, "badrum|NOUN": 8.44, "inbegripa|VERB": 8.44, "sovrum|NOUN": 8.44, "uppehålla|VERB": 8.44, "opassande|ADJ": 8.44, "hårddisk|NOUN": 8.43, "insamling|NOUN": 8.43, "oändligt|ADV": 8.43, "påminnelse|NOUN": 8.43, "marin|ADJ": 8.42, "opera|NOUN": 8.42, "aktieägare|NOUN": 8.41, "panel|NOUN": 8.41, "på något vis|ADV": 8.41, "inflytelserik|ADJ": 8.4, "polismyndighet|NOUN": 8.4, "vetenskapsman|NOUN": 8.4, "begåvad|ADJ": 8.4, "miljöfråga|NOUN": 8.39, "miste|PART": 8.39, "nicka|VERB": 8.39, "övervägande|ADJ": 8.39, "förtjänst|NOUN": 8.39, "inge|VERB": 8.39, "stolt|ADV": 8.39, "undergång|NOUN": 8.39, "ambitiös|ADJ": 8.38, "hebreisk|ADJ": 8.38, "växelkurs|NOUN": 8.38, "möda|NOUN": 8.37, "anklagad|ADJ": 8.37, "klassrum|NOUN": 8.36, "kontinuerlig|ADJ": 8.36, "si|ADV": 8.36, "entusiasm|NOUN": 8.35, "respons|NOUN": 8.35, "monster|NOUN": 8.34, "rån|NOUN": 8.34, "självkänsla|NOUN": 8.34, "sammanhållning|NOUN": 8.33, "sammanfalla|VERB": 8.32, "bara|SCONJ": 8.32, "intensivt|ADV": 8.32, "optimal|ADJ": 8.32, "suverän|ADJ": 8.32, "upp och ner|ADV": 8.32, "apotek|NOUN": 8.31, "hälla|VERB": 8.31, "käka|VERB": 8.31, "fäste|NOUN": 8.3, "hastigt|ADV": 8.3, "livslång|ADJ": 8.3, "svälta|VERB": 8.3, "välta|VERB": 8.3, "arbetsgivaravgift|NOUN": 8.29, "demon|NOUN": 8.29, "fastighetsskatt|NOUN": 8.29, "korridor|NOUN": 8.29, "stridsvagn|NOUN": 8.29, "tillvara|PART": 8.29, "vittnesmål|NOUN": 8.29, "ansvarsfull|ADJ": 8.28, "bagage|NOUN": 8.28, "evigt|ADV": 8.28, "koldioxidutsläpp|NOUN": 8.28, "fängsla|VERB": 8.27, "utflykt|NOUN": 8.27, "gratulera|VERB": 8.26, "studerande|NOUN": 8.26, "upprop|NOUN": 8.26, "utgåva|NOUN": 8.26, "vädja|VERB": 8.26, "finländsk|ADJ": 8.25, "morfar|NOUN": 8.25, "norrman|NOUN": 8.25, "skandinavisk|ADJ": 8.25, "tumme|NOUN": 8.25, "utslag|NOUN": 8.25, "familjemedlem|NOUN": 8.25, "lasta|VERB": 8.25, "ledarsida|NOUN": 8.25, "skräp|NOUN": 8.25, "smitta|VERB": 8.25, "påtala|VERB": 8.24, "stort|ADV": 8.24, "levnadsstandard|NOUN": 8.23, "palats|NOUN": 8.23, "tyska|NOUN": 8.23, "opinionsundersökning|NOUN": 8.22, "vetenskapligt|ADV": 8.22, "revidera|VERB": 8.22, "lovande|ADJ": 8.2, "orolighet|NOUN": 8.2, "brud|NOUN": 8.18, "tillvägagångssätt|NOUN": 8.18, "klistra|VERB": 8.18, "trams|NOUN": 8.18, "isär|PART": 8.17, "kärleksfull|ADJ": 8.17, "usch|INTJ": 8.16, "avslöjande|NOUN": 8.15, "beskatta|VERB": 8.15, "skrivbord|NOUN": 8.15, "utrikespolitisk|ADJ": 8.15, "vakta|VERB": 8.15, "arbetskamrat|NOUN": 8.14, "idiotisk|ADJ": 8.14, "spontant|ADV": 8.14, "tillställning|NOUN": 8.14, "tvärs|ADV": 8.14, "budgetår|NOUN": 8.13, "förtrycka|VERB": 8.13, "passande|ADJ": 8.13, "atom|NOUN": 8.12, "avta|VERB": 8.12, "chips|NOUN": 8.12, "markering|NOUN": 8.12, "tillåten|ADJ": 8.12, "öken|NOUN": 8.12, "sammanhängande|ADJ": 8.12, "fläck|NOUN": 8.11, "retorisk|ADJ": 8.11, "borgmästare|NOUN": 8.11, "förlorare|NOUN": 8.11, "melodi|NOUN": 8.11, "senat|NOUN": 8.11, "skarpt|ADV": 8.11, "sjöman|NOUN": 8.11, "bläddra|VERB": 8.1, "bärare|NOUN": 8.1, "gissning|NOUN": 8.1, "i onödan|ADV": 8.1, "stryk|NOUN": 8.1, "strålning|NOUN": 8.1, "terräng|NOUN": 8.1, "väva|VERB": 8.1, "skönt|ADV": 8.09, "spricka|VERB": 8.09, "äldreomsorg|NOUN": 8.09, "övertala|VERB": 8.09, "känslomässig|ADJ": 8.08, "feber|NOUN": 8.07, "härja|VERB": 8.07, "spelregel|NOUN": 8.07, "bekymrad|ADJ": 8.07, "annonsera|VERB": 8.06, "belastning|NOUN": 8.06, "flock|NOUN": 8.06, "inspektion|NOUN": 8.05, "laddning|NOUN": 8.05, "sammanslutning|NOUN": 8.05, "svek|NOUN": 8.05, "aska|NOUN": 8.04, "bekymra|VERB": 8.04, "finanspolitik|NOUN": 8.04, "godtycklig|ADJ": 8.04, "bluff|NOUN": 8.03, "distribuera|VERB": 8.03, "from|ADJ": 8.03, "förlopp|NOUN": 8.03, "nedläggning|NOUN": 8.03, "bestrida|VERB": 8.03, "huvudman|NOUN": 8.03, "ikapp|PART": 8.03, "empati|NOUN": 8.02, "sammansatt|ADJ": 8.01, "avlyssning|NOUN": 8.01, "dessförinnan|ADV": 8.01, "golf|NOUN": 8.01, "rasande|ADJ": 8.01, "reaktionär|ADJ": 8.01, "vifta|VERB": 8.0, "överklagande|NOUN": 8.0, "anor|NOUN": 7.99, "dominans|NOUN": 7.98, "lax|NOUN": 7.98, "organisering|NOUN": 7.98, "gift|NOUN": 7.97, "prostituerad|ADJ": 7.97, "återupprätta|VERB": 7.96, "hacka|VERB": 7.96, "medial|ADJ": 7.96, "entré|NOUN": 7.96, "farbror|NOUN": 7.96, "livlig|ADJ": 7.96, "packning|NOUN": 7.96, "essä|NOUN": 7.95, "magi|NOUN": 7.95, "självständigt|ADV": 7.95, "trötthet|NOUN": 7.95, "konsekvent|ADJ": 7.94, "rådgivning|NOUN": 7.94, "smälla|VERB": 7.94, "journalistisk|ADJ": 7.93, "officerare|NOUN": 7.93, "tjuv|NOUN": 7.93, "vidd|NOUN": 7.93, "belysning|NOUN": 7.92, "hänföra|VERB": 7.92, "nationalstat|NOUN": 7.92, "nedladdning|NOUN": 7.92, "växthuseffekt|NOUN": 7.92, "grotta|NOUN": 7.91, "matematisk|ADJ": 7.91, "ovanpå|ADP": 7.91, "pärla|NOUN": 7.91, "värk|NOUN": 7.91, "halvlek|NOUN": 7.9, "påtagligt|ADV": 7.9, "benägen|ADJ": 7.89, "recensera|VERB": 7.89, "diskriminera|VERB": 7.88, "pilot|NOUN": 7.88, "eftertanke|NOUN": 7.87, "fiktiv|ADJ": 7.87, "närliggande|ADJ": 7.87, "pålitlig|ADJ": 7.87, "korv|NOUN": 7.86, "reformera|VERB": 7.86, "pop|NOUN": 7.85, "fördubbla|VERB": 7.85, "militant|ADJ": 7.85, "sammantaget|ADV": 7.85, "tillkomst|NOUN": 7.85, "incident|NOUN": 7.84, "intill|ADV": 7.84, "underrättelse|NOUN": 7.84, "redigera|VERB": 7.83, "stadigt|ADV": 7.83, "baka|VERB": 7.82, "gud|INTJ": 7.82, "herregud|INTJ": 7.82, "observatör|NOUN": 7.82, "facit|NOUN": 7.82, "gruva|NOUN": 7.82, "obekväm|ADJ": 7.82, "fossil|ADJ": 7.81, "verkning|NOUN": 7.81, "kompromissa|VERB": 7.8, "konspirationsteori|NOUN": 7.8, "nacke|NOUN": 7.8, "svälja|VERB": 7.8, "tillstyrka|VERB": 7.8, "rättfärdighet|NOUN": 7.79, "adressat|NOUN": 7.79, "frågetecken|NOUN": 7.78, "image|NOUN": 7.78, "njutning|NOUN": 7.78, "utmärkt|ADV": 7.78, "isländsk|ADJ": 7.77, "skörda|VERB": 7.77, "såga|VERB": 7.77, "sökmotor|NOUN": 7.77, "drastiskt|ADV": 7.76, "dyrbar|ADJ": 7.76, "haka|VERB": 7.76, "knacka|VERB": 7.76, "offentlighet|NOUN": 7.76, "sekretess|NOUN": 7.76, "utkomma|VERB": 7.76, "indelning|NOUN": 7.75, "utomordentligt|ADV": 7.75, "olympisk|ADJ": 7.75, "skryta|VERB": 7.75, "ankomma|VERB": 7.74, "index|NOUN": 7.74, "umgänge|NOUN": 7.74, "välsignad|ADJ": 7.73, "avsky|VERB": 7.73, "förmoda|VERB": 7.73, "lyx|NOUN": 7.73, "skåp|NOUN": 7.72, "svamp|NOUN": 7.72, "uppehåll|NOUN": 7.72, "inbördes|ADJ": 7.71, "indikation|NOUN": 7.71, "jämlik|ADJ": 7.71, "staty|NOUN": 7.71, "uppförande|NOUN": 7.71, "överensstämmelse|NOUN": 7.71, "i grund och botten|ADV": 7.7, "puss|NOUN": 7.7, "spricka|NOUN": 7.7, "kemikalier|NOUN": 7.69, "konkurrenskraftig|ADJ": 7.69, "tankegång|NOUN": 7.69, "supporter|NOUN": 7.68, "symbolisk|ADJ": 7.68, "mervärde|NOUN": 7.68, "midsommar|NOUN": 7.68, "misstro|NOUN": 7.68, "fälla|NOUN": 7.67, "blues|NOUN": 7.66, "jury|NOUN": 7.66, "kör|NOUN": 7.66, "lyckligtvis|ADV": 7.66, "jordisk|ADJ": 7.65, "pumpa|VERB": 7.65, "harmoni|NOUN": 7.64, "trea|NOUN": 7.64, "avvägning|NOUN": 7.63, "markant|ADV": 7.62, "slopa|VERB": 7.62, "stål|NOUN": 7.62, "vinning|NOUN": 7.62, "främlingsfientlig|ADJ": 7.61, "mössa|NOUN": 7.61, "riksdagsman|NOUN": 7.61, "runtom|ADV": 7.61, "skikt|NOUN": 7.61, "avsevärd|ADJ": 7.61, "avvakta|VERB": 7.61, "dimma|NOUN": 7.61, "förundersökning|NOUN": 7.61, "huvudvärk|NOUN": 7.61, "ohälsa|NOUN": 7.61, "praktisera|VERB": 7.61, "rusta|VERB": 7.61, "subvention|NOUN": 7.61, "prisa|VERB": 7.61, "odemokratisk|ADJ": 7.6, "trilla|VERB": 7.6, "valfri|ADJ": 7.6, "mina|NOUN": 7.6, "ände|NOUN": 7.59, "hyresrätt|NOUN": 7.59, "härom|ADV": 7.59, "låga|NOUN": 7.59, "vital|ADJ": 7.59, "damm|NOUN": 7.3, "giftig|ADJ": 7.58, "pizza|NOUN": 7.58, "shopping|NOUN": 7.58, "färga|VERB": 7.58, "brygga|NOUN": 7.57, "kyckling|NOUN": 7.57, "löv|NOUN": 7.57, "specialist|NOUN": 7.57, "handlägga|VERB": 7.56, "hyckleri|NOUN": 7.56, "kännetecken|NOUN": 7.56, "överklass|NOUN": 7.56, "drivande|ADJ": 7.56, "arbetssätt|NOUN": 7.55, "hora|NOUN": 7.55, "nobelpris|NOUN": 7.55, "enkelhet|NOUN": 7.54, "förpliktelse|NOUN": 7.54, "larm|NOUN": 7.54, "lättnad|NOUN": 7.54, "predikan|NOUN": 7.54, "ammunition|NOUN": 7.53, "begär|NOUN": 7.53, "entydig|ADJ": 7.53, "missförstå|VERB": 7.53, "översvämning|NOUN": 7.53, "matcha|VERB": 7.53, "korrigera|VERB": 7.53, "försätta|VERB": 7.52, "frånvarande|ADJ": 7.51, "inblick|NOUN": 7.51, "ved|NOUN": 7.51, "mjukvara|NOUN": 7.5, "motpart|NOUN": 7.5, "riksdagsparti|NOUN": 7.5, "storskalig|ADJ": 7.5, "överflöd|NOUN": 7.5, "gröda|NOUN": 7.49, "jacka|NOUN": 7.49, "mottagande|NOUN": 7.49, "spårvagn|NOUN": 7.49, "återhämta|VERB": 7.49, "donera|VERB": 7.48, "sjukpenning|NOUN": 7.48, "bevarande|NOUN": 7.47, "bokhylla|NOUN": 7.47, "insida|NOUN": 7.47, "överraska|VERB": 7.47, "blöt|ADJ": 7.46, "relatera|VERB": 7.46, "underrättelsetjänst|NOUN": 7.46, "dynamik|NOUN": 7.46, "anmälning|NOUN": 7.45, "farhåga|NOUN": 7.45, "rovdjur|NOUN": 7.45, "tillsynsmyndighet|NOUN": 7.45, "adoptera|VERB": 7.45, "administrera|VERB": 7.44, "alltihop (vardagl. alltihopa)|PRON": 7.44, "dramatiskt|ADV": 7.44, "korkad|ADJ": 7.44, "marsch|NOUN": 7.44, "smäll|NOUN": 7.44, "less|ADJ": 7.43, "följande|ADJ": 7.42, "expedition|NOUN": 7.41, "heltäckande|ADJ": 7.41, "konvertera|VERB": 7.41, "i behov av|ADP": 7.4, "katastrofal|ADJ": 7.4, "näringsidkare|NOUN": 7.4, "otur|NOUN": 7.4, "flygning|NOUN": 7.39, "hierarki|NOUN": 7.39, "magasin|NOUN": 7.39, "plast|NOUN": 7.39, "stadig|ADJ": 7.39, "krävande|ADJ": 7.39, "täckt|ADJ": 7.39, "verifiera|VERB": 7.39, "blek|ADJ": 7.39, "förbjuden|ADJ": 7.39, "förnybar|ADJ": 7.39, "kyrkogård|NOUN": 7.39, "ovilja|NOUN": 7.39, "anarkist|NOUN": 7.38, "kartläggning|NOUN": 7.38, "krympa|VERB": 7.38, "skål|NOUN": 7.38, "underskatta|VERB": 7.38, "skifta|VERB": 7.37, "spänn|NOUN": 7.37, "auktion|NOUN": 7.36, "halka|VERB": 7.36, "kista|NOUN": 7.35, "sex|NOUN": 7.35, "vätska|NOUN": 7.34, "fascistisk|ADJ": 7.33, "hiss|NOUN": 7.33, "tå|NOUN": 7.33, "bestraffning|NOUN": 7.32, "bokstavligen|ADV": 7.32, "empirisk|ADJ": 7.32, "felaktigt|ADV": 7.32, "konfrontera|VERB": 7.32, "materia|NOUN": 7.32, "medborgerlig|ADJ": 7.32, "övergiven|ADJ": 7.32, "tillfredsställa|VERB": 7.32, "anmärkning|NOUN": 7.32, "nej|NOUN": 7.32, "skida|NOUN": 7.32, "förgäves|ADV": 7.31, "hiv|NOUN": 7.31, "kabel|NOUN": 7.31, "projektledare|NOUN": 7.31, "strikt|ADV": 7.31, "klinik|NOUN": 7.3, "råtta|NOUN": 7.3, "strömning|NOUN": 7.3, "kandidera|VERB": 7.29, "revolutionär|NOUN": 7.29, "ritning|NOUN": 7.29, "utmed|ADP": 7.29, "visdom|NOUN": 7.29, "uppfostra|VERB": 7.29, "lagändring|NOUN": 7.28, "så länge (som)|SCONJ": 7.28, "kulturarv|NOUN": 7.27, "nordlig|ADJ": 7.27, "plantera|VERB": 7.27, "chaufför|NOUN": 7.26, "inuti|ADP": 7.26, "förbruka|VERB": 7.25, "budgetproposition|NOUN": 7.25, "ceremoni|NOUN": 7.25, "uran|NOUN": 7.25, "aktualisera|VERB": 7.25, "barnfamilj|NOUN": 7.25, "population|NOUN": 7.25, "undanröja|VERB": 7.25, "utväg|NOUN": 7.25, "entreprenörskap|NOUN": 7.24, "godtagbar|ADJ": 7.24, "mardröm|NOUN": 7.24, "storebror|NOUN": 7.24, "isolera|VERB": 7.23, "kalas|NOUN": 7.23, "kopiering|NOUN": 7.23, "paroll|NOUN": 7.23, "shoppa|VERB": 7.23, "språkbruk|NOUN": 7.23, "diabetes|NOUN": 7.22, "fortlöpande|ADJ": 7.22, "klädsel|NOUN": 7.22, "svagt|ADV": 7.22, "ämbete|NOUN": 7.22, "historik|NOUN": 7.21, "intyg|NOUN": 7.21, "konversation|NOUN": 7.21, "växel|NOUN": 7.21, "byråkratisk|ADJ": 7.2, "etablering|NOUN": 7.2, "förnuftig|ADJ": 7.2, "hedra|VERB": 7.2, "omedveten|ADJ": 7.2, "stundtals|ADV": 7.2, "tjata|VERB": 7.2, "tjeckisk|ADJ": 7.2, "åtanke|NOUN": 7.2, "fördelaktig|ADJ": 7.19, "assistent|NOUN": 7.19, "läskig|ADJ": 7.19, "nationalekonomi|NOUN": 7.19, "återfå|VERB": 7.19, "övernaturlig|ADJ": 7.19, "elektricitet|NOUN": 7.18, "grovt|ADV": 7.18, "javisst (el. ja visst)|INTJ": 7.18, "beskylla|VERB": 7.18, "obegränsad|ADJ": 7.18, "anordning|NOUN": 7.18, "fluga|NOUN": 7.18, "förråd|NOUN": 7.18, "spänna|VERB": 7.18, "oönskad|ADJ": 7.18, "marschera|VERB": 7.17, "päls|NOUN": 7.17, "till vara|ADV": 7.17, "slant|NOUN": 7.16, "upprättande|NOUN": 7.16, "överdriva|VERB": 7.16, "reparera|VERB": 7.15, "central|NOUN": 7.15, "erövring|NOUN": 7.15, "justering|NOUN": 7.15, "nedanstående|ADJ": 7.15, "propagera|VERB": 7.15, "talesman|NOUN": 7.15, "uppträdande|NOUN": 7.15, "tandläkare|NOUN": 7.14, "utförande|NOUN": 7.14, "utgivare|NOUN": 7.14, "underordnad|ADJ": 7.14, "explosion|NOUN": 7.12, "fraktion|NOUN": 7.12, "renovera|VERB": 7.12, "snyggt|ADV": 7.12, "beröva|VERB": 7.11, "japan|NOUN": 7.11, "omvandling|NOUN": 7.11, "tillåtelse|NOUN": 7.11, "vidrig|ADJ": 7.11, "förmögen|ADJ": 7.11, "nedanför|ADP": 7.11, "oförmögen|ADJ": 7.11, "slösa|VERB": 7.11, "arbetsmarknadspolitik|NOUN": 7.1, "inkomstskatt|NOUN": 7.1, "skämta|VERB": 7.1, "underrätta|VERB": 7.1, "världslig|ADJ": 7.1, "cigarett|NOUN": 7.09, "hälsosam|ADJ": 7.09, "skalle|NOUN": 7.09, "spädbarn|NOUN": 7.09, "domslut|NOUN": 7.08, "dyrka|VERB": 7.08, "utmärkelse|NOUN": 7.08, "katalog|NOUN": 7.07, "bredband|NOUN": 7.07, "kemi|NOUN": 7.07, "foster|NOUN": 7.06, "tillfällighet|NOUN": 7.06, "enastående|ADJ": 7.05, "rökning|NOUN": 7.05, "trots|NOUN": 7.05, "muta|NOUN": 7.04, "motgång|NOUN": 7.04, "människosyn|NOUN": 7.04, "omvända|VERB": 7.04, "sammanbrott|NOUN": 7.04, "auktoritär|ADJ": 7.03, "bebis|NOUN": 7.03, "fat|NOUN": 7.03, "hunger|NOUN": 7.03, "metafor|NOUN": 7.03, "understödja|VERB": 7.03, "anamma|VERB": 7.03, "arrestera|VERB": 7.03, "barriär|NOUN": 7.02, "best|NOUN": 7.02, "fästning|NOUN": 7.02, "immateriell|ADJ": 7.02, "vansinne|NOUN": 7.02, "involvera|VERB": 7.02, "hopplös|ADJ": 7.01, "införliva|VERB": 7.01, "tacksamhet|NOUN": 7.01, "återkalla|VERB": 7.01, "jämnt|ADJ": 7.0, "extremist|NOUN": 7.0, "civilbefolkning|NOUN": 6.99, "förtvivlan|NOUN": 6.99, "löntagare|NOUN": 6.99, "åratal|NOUN": 6.99, "överträffa|VERB": 6.99, "flitig|ADJ": 6.99, "härleda|VERB": 6.98, "greve|NOUN": 6.98, "internt|ADV": 6.98, "soppa|NOUN": 6.98, "tvivelaktig|ADJ": 6.98, "ändamålsenlig|ADJ": 6.98, "byråkrat|NOUN": 6.97, "lagstiftande|ADJ": 6.97, "civiliserad|ADJ": 6.97, "fjäll|NOUN": 6.97, "knäcka|VERB": 6.97, "likgiltig|ADJ": 6.97, "nationalist|NOUN": 6.97, "offensiv|ADJ": 6.97, "socialbidrag|NOUN": 6.97, "befästa|VERB": 6.96, "väninna|NOUN": 6.96, "blixt|NOUN": 6.96, "bevisligen|ADV": 6.96, "fräsch|ADJ": 6.96, "ivrig|ADJ": 6.96, "mus|NOUN": 6.96, "tillkännagivande|NOUN": 6.96, "lojal|ADJ": 6.95, "småföretag|NOUN": 6.95, "terapi|NOUN": 6.95, "undanta|VERB": 6.95, "frekvens|NOUN": 6.94, "givande|ADJ": 6.94, "i ljuset av|ADP": 6.94, "komisk|ADJ": 6.94, "kostnadsfri|ADJ": 6.94, "uniform|NOUN": 6.94, "utfrågning|NOUN": 6.94, "godhet|NOUN": 6.93, "tysta|VERB": 6.93, "bombning|NOUN": 6.92, "engelskspråkig|ADJ": 6.92, "beslag|NOUN": 6.91, "vapenvila|NOUN": 6.91, "buller|NOUN": 6.9, "intervention|NOUN": 6.9, "lagring|NOUN": 6.9, "utbyta|VERB": 6.9, "svin|NOUN": 6.9, "lagom|ADJ": 6.89, "doktrin|NOUN": 6.89, "klick|NOUN": 6.89, "stämpla|VERB": 6.89, "uppfostran|NOUN": 6.89, "bilateral|ADJ": 6.88, "bostadsrätt|NOUN": 6.88, "iakttagelse|NOUN": 6.88, "på sistone|ADV": 6.88, "påskynda|VERB": 6.88, "sponsra|VERB": 6.88, "avbrott|NOUN": 6.87, "bestånd|NOUN": 6.87, "hantverkare|NOUN": 6.87, "sjukskrivning|NOUN": 6.87, "slakta|VERB": 6.87, "uppröra|VERB": 6.87, "besittning|NOUN": 6.86, "fasa|NOUN": 6.86, "konfrontation|NOUN": 6.86, "trådlös|ADJ": 6.86, "pub|NOUN": 6.85, "biverkning|NOUN": 6.85, "dragning|NOUN": 6.85, "logiskt|ADV": 6.85, "österut|ADV": 6.85, "deckare|NOUN": 6.84, "dåtid|NOUN": 6.84, "cynisk|ADJ": 6.83, "poetisk|ADJ": 6.83, "kostsam|ADJ": 6.82, "misslyckad|ADJ": 6.82, "prioritet|NOUN": 6.82, "fascist|NOUN": 6.82, "frestelse|NOUN": 6.82, "trösta|VERB": 6.82, "uppriktigt|ADV": 6.82, "världsekonomi|NOUN": 6.82, "summera|VERB": 6.82, "fängelsestraff|NOUN": 6.81, "invigning|NOUN": 6.81, "revisor|NOUN": 6.81, "samisk|ADJ": 6.81, "så snart som|ADV": 6.81, "underminera|VERB": 6.81, "medgivande|NOUN": 6.8, "tvätt|NOUN": 6.8, "guvernör|NOUN": 6.8, "adekvat|ADJ": 6.79, "brottas|VERB": 6.79, "hantverk|NOUN": 6.79, "minus|ADV": 6.79, "fullborda|VERB": 6.79, "latinsk|ADJ": 6.78, "stabilisera|VERB": 6.78, "kvantitet|NOUN": 6.78, "huvudroll|NOUN": 6.77, "hög|NOUN": 6.77, "knepig|ADJ": 6.77, "överblick|NOUN": 6.77, "berömma|VERB": 6.77, "räckvidd|NOUN": 6.76, "utifrån|ADV": 6.76, "västlig|ADJ": 6.76, "skicklighet|NOUN": 6.75, "bestraffa|VERB": 6.75, "spik|NOUN": 6.75, "akademiker|NOUN": 6.75, "författarskap|NOUN": 6.75, "närvara|VERB": 6.75, "sola|VERB": 6.74, "association|NOUN": 6.74, "exil|NOUN": 6.74, "förbehåll|NOUN": 6.74, "hämma|VERB": 6.74, "nominera|VERB": 6.74, "viska|VERB": 6.74, "koalition|NOUN": 6.73, "spektakulär|ADJ": 6.73, "teoretiskt|ADV": 6.73, "handfull|NOUN": 6.72, "ugn|NOUN": 6.72, "geografi|NOUN": 6.72, "meditation|NOUN": 6.72, "betoning|NOUN": 6.71, "brevlåda|NOUN": 6.71, "förfoga|VERB": 6.71, "heja|VERB": 6.71, "ironisk|ADJ": 6.71, "skrivare|NOUN": 6.71, "valdeltagande|NOUN": 6.71, "lamm|NOUN": 6.7, "berika|VERB": 6.7, "brytning|NOUN": 6.7, "flyktingpolitik|NOUN": 6.7, "porr|NOUN": 6.7, "flöda|VERB": 6.69, "revolt|NOUN": 6.69, "snällt|ADV": 6.69, "vika|ADV": 6.69, "ekosystem|NOUN": 6.68, "heterosexuell|ADJ": 6.68, "kolumn|NOUN": 6.68, "lyssnare|NOUN": 6.68, "möjligt|ADV": 6.68, "utebli|VERB": 6.68, "underkasta|VERB": 6.68, "salong|NOUN": 6.68, "sjöfart|NOUN": 6.68, "tapet|NOUN": 6.68, "bråttom|ADV": 6.67, "kraftverk|NOUN": 6.67, "spotta|VERB": 6.67, "duscha|VERB": 6.66, "attrahera|VERB": 6.66, "måste|NOUN": 6.66, "ovannämnd|ADJ": 6.66, "tänkare|NOUN": 6.66, "morot|NOUN": 6.65, "censurera|VERB": 6.65, "lagtext|NOUN": 6.65, "lindra|VERB": 6.65, "vilse|ADV": 6.65, "förenkling|NOUN": 6.64, "tolerera|VERB": 6.64, "löst|ADV": 6.64, "sankt (förk. s:t)|ADJ": 6.64, "överflödig|ADJ": 6.64, "omnämna|VERB": 6.63, "pund|NOUN": 6.63, "slöseri|NOUN": 6.63, "formel|NOUN": 6.62, "drink|NOUN": 6.62, "förväntan|NOUN": 6.62, "lunga|NOUN": 6.62, "vårdcentral|NOUN": 6.62, "ödmjukhet|NOUN": 6.62, "överdrift|NOUN": 6.62, "häpnadsväckande|ADJ": 6.61, "urskilja|VERB": 6.61, "frigörelse|NOUN": 6.61, "monetär|ADJ": 6.61, "tobak|NOUN": 6.61, "tråkigt|ADV": 6.61, "förordna|VERB": 6.61, "femma|NOUN": 6.61, "livslängd|NOUN": 6.61, "sval|ADJ": 6.61, "telefonnummer|NOUN": 6.61, "analytiker|NOUN": 6.6, "avspegla|VERB": 6.6, "psykiatrisk|ADJ": 6.6, "rebell|NOUN": 6.6, "droppa|VERB": 6.59, "tugga|VERB": 6.59, "kval|NOUN": 6.59, "läroplan|NOUN": 6.59, "psalm|NOUN": 6.59, "sårbar|ADJ": 6.59, "kår|NOUN": 6.58, "luthersk|ADJ": 6.58, "stel|ADJ": 6.58, "tydliggöra|VERB": 6.58, "barnslig|ADJ": 6.57, "betraktelse|NOUN": 6.57, "fortgå|VERB": 6.57, "optimistisk|ADJ": 6.57, "tillfredsställelse|NOUN": 6.57, "välmående|ADJ": 6.57, "applicera|VERB": 6.56, "förkortning|NOUN": 6.56, "jämställa|VERB": 6.56, "runt omkring|ADV": 6.56, "välsigna|VERB": 6.56, "donation|NOUN": 6.56, "laddad|ADJ": 6.56, "monument|NOUN": 6.55, "blomma|VERB": 6.55, "hona|NOUN": 6.55, "prick|NOUN": 6.55, "humanistisk|ADJ": 6.54, "intressent|NOUN": 6.54, "parameter|NOUN": 6.54, "sopa|VERB": 6.54, "streck|NOUN": 6.54, "ikon|NOUN": 6.54, "insekt|NOUN": 6.54, "dotterbolag|NOUN": 6.53, "irakier|NOUN": 6.53, "istid|NOUN": 6.53, "till slut|ADV": 6.53, "försening|NOUN": 6.53, "färja|NOUN": 6.53, "förståelig|ADJ": 6.53, "prenumerera|VERB": 6.53, "ansluten|ADJ": 6.53, "romantik|NOUN": 6.53, "bisarr|ADJ": 6.52, "förfalla|VERB": 6.52, "lås|NOUN": 6.52, "principiellt|ADV": 6.52, "samförstånd|NOUN": 6.52, "jazz|NOUN": 6.52, "ritual|NOUN": 6.52, "segel|NOUN": 6.51, "exotisk|ADJ": 6.51, "informationssamhälle|NOUN": 6.51, "lukt|NOUN": 6.51, "skrapa|VERB": 6.51, "uppgradera|VERB": 6.51, "mäklare|NOUN": 6.51, "reservera|VERB": 6.51, "bur|NOUN": 6.5, "snöa|VERB": 6.5, "anteckna|VERB": 6.5, "box|NOUN": 6.5, "korsning|NOUN": 6.5, "legitimera|VERB": 6.5, "förfärlig|ADJ": 6.49, "förvånansvärt|ADV": 6.49, "kretsa|VERB": 6.49, "implementera|VERB": 6.48, "alster|NOUN": 6.48, "energikälla|NOUN": 6.48, "livsfarlig|ADJ": 6.48, "livskvalitet|NOUN": 6.48, "måttlig|ADJ": 6.48, "tryggt|ADV": 6.48, "bäck|NOUN": 6.47, "förtal|NOUN": 6.47, "förutsägbar|ADJ": 6.47, "intensifiera|VERB": 6.47, "naturresurs|NOUN": 6.47, "otänkbar|ADJ": 6.47, "varsel|NOUN": 6.47, "tillbehör|NOUN": 6.47, "betong|NOUN": 6.46, "nybörjare|NOUN": 6.46, "ruin|NOUN": 6.46, "sortiment|NOUN": 6.46, "nyans|NOUN": 6.46, "uppbära|VERB": 6.46, "arkeologisk|ADJ": 6.46, "okunnighet|NOUN": 6.46, "anseende|NOUN": 6.46, "förbannelse|NOUN": 6.46, "jubla|VERB": 6.46, "lejon|NOUN": 6.46, "session|NOUN": 6.46, "effektivisera|VERB": 6.45, "hotfull|ADJ": 6.45, "miljöpolitik|NOUN": 6.45, "storföretag|NOUN": 6.45, "suveränitet|NOUN": 6.45, "utanför|ADV": 6.45, "landshövding|NOUN": 6.45, "statsbidrag|NOUN": 6.44, "storslagen|ADJ": 6.44, "separera|VERB": 6.43, "firande|NOUN": 6.43, "hyllning|NOUN": 6.43, "oljepris|NOUN": 6.43, "biologi|NOUN": 6.42, "rimligtvis|ADV": 6.42, "arbetarparti|NOUN": 6.41, "beskåda|VERB": 6.41, "briljant|ADJ": 6.41, "lott|NOUN": 6.41, "kidnappa|VERB": 6.41, "girighet|NOUN": 6.4, "härröra|VERB": 6.4, "på sätt och vis|ADV": 6.4, "framlägga|VERB": 6.4, "förorsaka|VERB": 6.4, "häck|NOUN": 6.4, "hemvist|NOUN": 6.4, "andetag|NOUN": 6.39, "berusad|ADJ": 6.39, "tortera|VERB": 6.39, "kanadensisk|ADJ": 6.39, "protestantisk|ADJ": 6.39, "läktare|NOUN": 6.39, "marxist|NOUN": 6.39, "peta|VERB": 6.39, "sakkunnig|ADJ": 6.39, "svängning|NOUN": 6.39, "tanka|VERB": 6.39, "sympatisk|ADJ": 6.39, "översikt|NOUN": 6.39, "midnatt|NOUN": 6.38, "amatör|NOUN": 6.38, "befalla|VERB": 6.37, "handledare|NOUN": 6.37, "bostadsmarknad|NOUN": 6.37, "klappa|VERB": 6.37, "media|NOUN": 6.37, "när som helst|ADV": 6.37, "pil|NOUN": 6.37, "rättsstat|NOUN": 6.37, "röra|NOUN": 6.37, "vålla|VERB": 6.36, "blygsam|ADJ": 6.36, "exponering|NOUN": 6.36, "närområde|NOUN": 6.36, "otrogen|ADJ": 6.36, "varva|VERB": 6.36, "regent|NOUN": 6.35, "bunt|NOUN": 6.35, "fostra|VERB": 6.35, "funktionell|ADJ": 6.35, "klinisk|ADJ": 6.35, "värdegrund|NOUN": 6.35, "förutsäga|VERB": 6.35, "begrunda|VERB": 6.34, "tennis|NOUN": 6.34, "destination|NOUN": 6.34, "taktisk|ADJ": 6.34, "österrikisk|ADJ": 6.34, "manifestera|VERB": 6.34, "förakta|VERB": 6.33, "invandringspolitik|NOUN": 6.33, "utbrista|VERB": 6.33, "aids|NOUN": 6.33, "bekanta|VERB": 6.33, "utövare|NOUN": 6.32, "angå|VERB": 6.32, "förlossning|NOUN": 6.32, "återgång|NOUN": 6.32, "procedur|NOUN": 6.32, "äventyra|VERB": 6.32, "rep|NOUN": 6.31, "sväva|VERB": 6.31, "diet|NOUN": 6.31, "filter|NOUN": 6.31, "gratis|ADJ": 6.31, "legendarisk|ADJ": 6.31, "plagg|NOUN": 6.31, "impuls|NOUN": 6.3, "parkering|NOUN": 6.3, "beståndsdel|NOUN": 6.3, "brottslig|ADJ": 6.3, "årstid|NOUN": 6.3, "underlåta|VERB": 6.29, "episod|NOUN": 6.28, "kock|NOUN": 6.28, "affärsman|NOUN": 6.28, "högkonjunktur|NOUN": 6.28, "lur|NOUN": 6.28, "nu|NOUN": 6.28, "opinionsbildning|NOUN": 6.28, "premiss|NOUN": 6.28, "insistera|VERB": 6.28, "grafik|NOUN": 6.27, "munk|NOUN": 6.27, "skörd|NOUN": 6.27, "dräkt|NOUN": 6.27, "galenskap|NOUN": 6.27, "franska|NOUN": 6.27, "pistol|NOUN": 6.27, "pyssla|VERB": 6.27, "urholka|VERB": 6.27, "galning|NOUN": 6.26, "hugg|NOUN": 6.26, "preferens|NOUN": 6.26, "uppslag|NOUN": 6.26, "exploatera|VERB": 6.26, "förväxla|VERB": 6.26, "tomat|NOUN": 6.26, "ocean|NOUN": 6.26, "cyklist|NOUN": 6.25, "näve|NOUN": 6.25, "omstrukturering|NOUN": 6.25, "restriktiv|ADJ": 6.25, "skina|VERB": 6.25, "skulptur|NOUN": 6.25, "ättling|NOUN": 6.25, "helgon|NOUN": 6.25, "utstå|VERB": 6.25, "envisas|VERB": 6.25, "pedagogik|NOUN": 6.25, "postning|NOUN": 6.25, "trygga|VERB": 6.25, "uppmärksam|ADJ": 6.25, "bädda|VERB": 6.24, "fuktig|ADJ": 6.24, "fundament|NOUN": 6.24, "reformation|NOUN": 6.24, "grilla|VERB": 6.23, "italienare|NOUN": 6.23, "famn|NOUN": 6.23, "genomgripande|ADJ": 6.23, "skägg|NOUN": 6.23, "slappna|VERB": 6.23, "medalj|NOUN": 6.23, "expansiv|ADJ": 6.22, "matlagning|NOUN": 6.22, "rytm|NOUN": 6.22, "elefant|NOUN": 6.22, "patetisk|ADJ": 6.22, "batteri|NOUN": 6.22, "tippa|VERB": 6.22, "ambulans|NOUN": 6.21, "bearbetning|NOUN": 6.21, "huvudkontor|NOUN": 6.21, "precisera|VERB": 6.21, "folkmassa|NOUN": 6.21, "ohållbar|ADJ": 6.21, "revision|NOUN": 6.21, "såra|VERB": 6.21, "mix|NOUN": 6.21, "vy|NOUN": 6.21, "diplomat|NOUN": 6.2, "affisch|NOUN": 6.2, "associera|VERB": 6.2, "kalkyl|NOUN": 6.2, "konstgjord|ADJ": 6.2, "polack|NOUN": 6.2, "renovering|NOUN": 6.2, "maffia|NOUN": 6.19, "snickare|NOUN": 6.19, "teolog|NOUN": 6.19, "väster om|ADP": 6.19, "kontinuitet|NOUN": 6.19, "marginell|ADJ": 6.19, "ojämn|ADJ": 6.19, "skoja|VERB": 6.18, "tangentbord|NOUN": 6.18, "migration|NOUN": 6.18, "säck|NOUN": 6.18, "körning|NOUN": 6.18, "blond|ADJ": 6.18, "dygd|NOUN": 6.18, "förorening|NOUN": 6.18, "svenskspråkig|ADJ": 6.18, "lera|NOUN": 6.18, "befattning|NOUN": 6.17, "föredöme|NOUN": 6.17, "genetiskt|ADV": 6.17, "sucka|VERB": 6.17, "framhäva|VERB": 6.17, "laboratorium|NOUN": 6.17, "strypa|VERB": 6.17, "kroppslig|ADJ": 6.16, "pool|NOUN": 6.16, "sionism|NOUN": 6.16, "uttag|NOUN": 6.16, "begynnelse|NOUN": 6.15, "likartad|ADJ": 6.15, "slakt|NOUN": 6.15, "naturvetenskap|NOUN": 6.14, "premie|NOUN": 6.14, "snus|NOUN": 6.14, "tillgå|VERB": 6.14, "vadå|INTJ": 6.14, "valresultat|NOUN": 6.14, "västerut|ADV": 6.14, "diamant|NOUN": 6.14, "kulle|NOUN": 6.14, "avlyssna|VERB": 6.13, "bärbar|ADJ": 6.13, "förkylning|NOUN": 6.13, "piano|NOUN": 6.13, "plåga|NOUN": 6.13, "signalera|VERB": 6.13, "snubbe|NOUN": 6.13, "eftergift|NOUN": 6.13, "major|NOUN": 6.13, "veterinär|NOUN": 6.13, "utopi|NOUN": 6.12, "författa|VERB": 6.12, "gräsmatta|NOUN": 6.12, "bifoga|VERB": 6.11, "parkera|VERB": 6.11, "fastland|NOUN": 6.11, "mentalitet|NOUN": 6.11, "slagfält|NOUN": 6.11, "stimulans|NOUN": 6.11, "proffs|NOUN": 6.11, "ekvation|NOUN": 6.1, "repris|NOUN": 6.1, "rådgivande|ADJ": 6.1, "vinnande|ADJ": 6.1, "diskret|ADJ": 6.09, "befallning|NOUN": 6.09, "pipa|NOUN": 6.09, "kjol|NOUN": 6.08, "bubbla|NOUN": 6.08, "mirakel|NOUN": 6.08, "hednisk|ADJ": 6.07, "lök|NOUN": 6.07, "infektion|NOUN": 6.06, "integrering|NOUN": 6.06, "uträtta|VERB": 6.06, "älskling|NOUN": 6.06, "pedagog|NOUN": 6.06, "kvalitativ|ADJ": 6.05, "motorcykel|NOUN": 6.05, "styrelseledamot|NOUN": 6.04, "tvärt|ADV": 6.04, "domän|NOUN": 6.04, "subjekt|NOUN": 6.03, "fana|NOUN": 6.03, "fax|NOUN": 0.79, "belasta|VERB": 6.02, "föreläsare|NOUN": 6.01, "lagstiftare|NOUN": 6.01, "högkvarter|NOUN": 6.0, "fascinera|VERB": 5.99, "fånig|ADJ": 5.99, "administratör|NOUN": 5.99, "förälskad|ADJ": 5.98, "gagna|VERB": 5.98, "modifiera|VERB": 5.98, "realisera|VERB": 5.98, "samlag|NOUN": 5.98, "skymta|VERB": 5.98, "utbredning|NOUN": 5.98, "utkant|NOUN": 5.97, "envis|ADJ": 5.97, "syndare|NOUN": 5.96, "paradox|NOUN": 5.96, "bräda|NOUN": 5.96, "ordbok|NOUN": 5.96, "översättare|NOUN": 5.96, "avkomma|NOUN": 5.95, "avlägga|VERB": 5.95, "utnämning|NOUN": 5.95, "riddare|NOUN": 5.95, "handikapp|NOUN": 5.94, "myra|NOUN": 5.94, "hop|NOUN": 5.93, "föreläsa|VERB": 5.93, "besläktad|ADJ": 5.92, "halvö|NOUN": 5.92, "sammanslagning|NOUN": 5.92, "yngling|NOUN": 5.92, "klassificera|VERB": 5.91, "spruta|VERB": 5.91, "spärra|VERB": 5.91, "biograf|NOUN": 5.9, "klan|NOUN": 5.9, "löpning|NOUN": 5.9, "profit|NOUN": 5.9, "hållbarhet|NOUN": 5.89, "foder|NOUN": 5.89, "framsida|NOUN": 5.89, "solidarisk|ADJ": 5.89, "tallrik|NOUN": 5.89, "nominering|NOUN": 5.88, "handbok|NOUN": 5.88, "debut|NOUN": 5.87, "försiktighet|NOUN": 5.87, "groda|NOUN": 5.87, "hobby|NOUN": 5.86, "bidragande|ADJ": 5.85, "blomstra|VERB": 5.85, "välbefinnande|NOUN": 5.85, "deg|NOUN": 5.84, "demo|NOUN": 5.84, "fiskare|NOUN": 5.84, "ryggsäck|NOUN": 5.84, "behaga|VERB": 5.84, "ekumenisk|ADJ": 5.84, "partikel|NOUN": 5.84, "svettig|ADJ": 5.84, "tårta|NOUN": 5.84, "utsida|NOUN": 5.84, "drunkna|VERB": 5.83, "kognitiv|ADJ": 5.83, "prägel|NOUN": 5.83, "klang|NOUN": 5.83, "pc|NOUN": 5.83, "faktura|NOUN": 5.82, "oroväckande|ADJ": 5.82, "broschyr|NOUN": 5.82, "mästerskap|NOUN": 5.82, "terror|NOUN": 5.82, "duk|NOUN": 5.8, "expertis|NOUN": 5.8, "jungfru|NOUN": 5.8, "utgivning|NOUN": 5.78, "avundsjuka|NOUN": 5.77, "multinationell|ADJ": 5.77, "vett|NOUN": 5.76, "insättning|NOUN": 5.75, "statisk|ADJ": 5.75, "stavning|NOUN": 5.75, "steka|VERB": 5.74, "bedra|VERB": 5.74, "förvandling|NOUN": 5.74, "snäv|ADJ": 5.73, "läka|VERB": 5.72, "nagel|NOUN": 5.72, "utdragen|ADJ": 5.72, "överordnad|ADJ": 5.71, "tillbe|VERB": 5.7, "avsändare|NOUN": 5.7, "beklaglig|ADJ": 5.7, "sköld|NOUN": 5.69, "syre|NOUN": 5.69, "bubbla|VERB": 5.68, "kväva|VERB": 5.68, "motstå|VERB": 5.68, "väktare|NOUN": 5.68, "express|NOUN": 5.67, "häxa|NOUN": 5.67, "irritera|VERB": 5.66, "lärobok|NOUN": 5.66, "nerv|NOUN": 5.65, "pendla|VERB": 5.65, "trakassera|VERB": 5.65, "förvaring|NOUN": 5.64, "oskuld|NOUN": 5.64, "sydlig|ADJ": 5.64, "gudinna|NOUN": 5.64, "sponsor|NOUN": 5.64, "bekantskap|NOUN": 5.63, "skoj|ADJ": 5.63, "filial|NOUN": 5.62, "kvalifikation|NOUN": 5.62, "ratificera|VERB": 5.62, "spis|NOUN": 5.62, "strumpa|NOUN": 5.62, "hetta|NOUN": 5.61, "kyssa|VERB": 5.61, "sekundär|ADJ": 5.61, "utmanande|ADJ": 5.61, "avbilda|VERB": 5.61, "segling|NOUN": 5.61, "drastisk|ADJ": 5.6, "korg|NOUN": 5.6, "avsiktligt|ADV": 5.59, "tystna|VERB": 5.59, "underjordisk|ADJ": 5.59, "entusiastisk|ADJ": 5.58, "talarstol|NOUN": 5.58, "omöjlighet|NOUN": 5.57, "kriga|VERB": 5.57, "kylskåp|NOUN": 5.57, "skoj|NOUN": 5.57, "omkomma|VERB": 5.56, "territoriell|ADJ": 5.56, "provisorisk|ADJ": 5.55, "tablett|NOUN": 5.55, "galax|NOUN": 5.55, "sallad|NOUN": 5.55, "berömd|ADJ": 5.54, "hjälm|NOUN": 5.54, "teknologisk|ADJ": 5.54, "försumma|VERB": 5.53, "föråldrad|ADJ": 5.53, "komplexitet|NOUN": 5.53, "kronisk|ADJ": 5.53, "geni|NOUN": 5.53, "kvadratmeter|NOUN": 5.52, "tillfoga|VERB": 5.52, "upprepning|NOUN": 5.51, "cirkulera|VERB": 5.5, "kvantitativ|ADJ": 5.5, "kvot|NOUN": 5.5, "hallå|INTJ": 5.47, "tröskel|NOUN": 5.47, "syndrom|NOUN": 5.47, "tvilling|NOUN": 5.47, "modernisera|VERB": 5.46, "stämpel|NOUN": 5.46, "autonomi|NOUN": 5.46, "mjöl|NOUN": 5.46, "vägledande|ADJ": 5.46, "slagsmål|NOUN": 5.45, "semifinal|NOUN": 5.45, "diktera|VERB": 5.44, "lärorik|ADJ": 5.44, "samarbetspartner|NOUN": 5.44, "envar|PRON": 5.44, "bokhandel|NOUN": 5.43, "dunkel|ADJ": 5.43, "reparation|NOUN": 5.43, "docka|NOUN": 5.43, "obehag|NOUN": 5.43, "originell|ADJ": 5.43, "galleri|NOUN": 5.42, "ökänd|ADJ": 5.42, "mottagning|NOUN": 5.42, "intensitet|NOUN": 5.41, "modernisering|NOUN": 5.41, "visuell|ADJ": 5.4, "kommentator|NOUN": 5.4, "beskydd|NOUN": 5.4, "döv|ADJ": 5.39, "knäppa|VERB": 5.39, "grundlig|ADJ": 5.39, "husdjur|NOUN": 5.39, "halvvägs|ADV": 5.37, "tomhet|NOUN": 5.37, "ansats|NOUN": 5.36, "iskall|ADJ": 5.36, "ofattbar|ADJ": 5.36, "tiger|NOUN": 5.36, "applikation|NOUN": 5.36, "självstyre|NOUN": 5.36, "mästerverk|NOUN": 5.35, "svett|NOUN": 5.35, "studsa|VERB": 5.34, "optimism|NOUN": 5.33, "uppgradering|NOUN": 5.33, "befordra|VERB": 5.33, "intyga|VERB": 5.33, "vinka|VERB": 5.33, "motsägelse|NOUN": 5.32, "martyr|NOUN": 5.32, "satellit|NOUN": 5.32, "uppriktig|ADJ": 5.31, "bedrift|NOUN": 5.3, "förvaltare|NOUN": 5.3, "biträdande|ADJ": 5.3, "segrare|NOUN": 5.29, "dumpa|VERB": 5.28, "övervikt|NOUN": 5.28, "kollapsa|VERB": 5.27, "städning|NOUN": 5.27, "borra|VERB": 5.26, "nyfödd|ADJ": 5.26, "smink|NOUN": 5.26, "parentes|NOUN": 5.25, "infödd|ADJ": 5.25, "irritation|NOUN": 5.25, "rutten|ADJ": 5.25, "fakultet|NOUN": 5.25, "skiss|NOUN": 5.25, "rand|NOUN": 5.25, "festa|VERB": 5.24, "frekvent|ADJ": 5.24, "prestanda|NOUN": 5.24, "djärv|ADJ": 5.24, "omtyckt|ADJ": 5.24, "skrik|NOUN": 5.23, "förtvivlad|ADJ": 5.23, "uttrycklig|ADJ": 5.23, "signera|VERB": 5.22, "experimentera|VERB": 5.21, "födsel|NOUN": 5.21, "ombyggnad|NOUN": 5.2, "avgrund|NOUN": 5.19, "kapell|NOUN": 5.19, "planta|NOUN": 5.19, "våt|ADJ": 5.18, "fångenskap|NOUN": 5.18, "korrekthet|NOUN": 5.18, "variabel|NOUN": 5.18, "formulär|NOUN": 5.18, "gap|NOUN": 5.18, "manifest|NOUN": 5.18, "handlare|NOUN": 5.17, "mobilisering|NOUN": 5.17, "återförsäljare|NOUN": 5.17, "fördjupning|NOUN": 5.16, "räv|NOUN": 5.16, "anvisa|VERB": 5.16, "definitiv|ADJ": 5.16, "misstänksam|ADJ": 5.16, "intervall|NOUN": 5.15, "gryta|NOUN": 5.15, "återvinna|VERB": 5.15, "frakta|VERB": 5.14, "gumma|NOUN": 5.14, "ojämlikhet|NOUN": 5.14, "krut|NOUN": 5.14, "precision|NOUN": 5.14, "anslå|VERB": 5.13, "orealistisk|ADJ": 5.13, "copyright|NOUN": 5.13, "företräde|NOUN": 5.13, "minimum|NOUN": 5.13, "skolgång|NOUN": 5.12, "giltighet|NOUN": 5.11, "anknyta|VERB": 5.11, "avskeda|VERB": 5.11, "barmhärtighet|NOUN": 5.11, "gevär|NOUN": 5.11, "visum|NOUN": 5.11, "analytisk|ADJ": 5.1, "intrig|NOUN": 5.1, "förkorta|VERB": 5.09, "påträffa|VERB": 5.09, "skådespel|NOUN": 5.09, "avtryck|NOUN": 5.07, "disponera|VERB": 5.07, "knuffa|VERB": 5.07, "vägran|NOUN": 5.07, "charm|NOUN": 5.05, "uthärda|VERB": 5.05, "högtidlig|ADJ": 5.05, "komplikation|NOUN": 5.05, "delegat|NOUN": 5.04, "socialförsäkring|NOUN": 5.04, "öm|ADJ": 5.04, "bälte|NOUN": 5.03, "privatisera|VERB": 5.03, "lillebror|NOUN": 5.03, "smuts|NOUN": 5.03, "kudde|NOUN": 5.02, "slätt|NOUN": 5.02, "kondom|NOUN": 5.01, "tank|NOUN": 5.01, "bråkdel|NOUN": 5.01, "ögonbryn|NOUN": 5.01, "undkomma|VERB": 4.99, "hejdå (el. hej då)|INTJ": 4.99, "spannmål|NOUN": 4.97, "uttal|NOUN": 4.97, "kompositör|NOUN": 4.97, "korn|NOUN": 4.97, "täckning|NOUN": 4.97, "anstalt|NOUN": 4.96, "förmedling|NOUN": 4.96, "deprimerad|ADJ": 4.95, "sammankomst|NOUN": 4.95, "vänligen|ADV": 4.95, "grymhet|NOUN": 4.94, "nykter|ADJ": 4.93, "solid|ADJ": 4.92, "idealisk|ADJ": 4.92, "pyramid|NOUN": 4.92, "stövel|NOUN": 4.92, "gråt|NOUN": 4.9, "täcke|NOUN": 4.9, "blinka|VERB": 4.9, "gränd|NOUN": 4.9, "otillåten|ADJ": 4.9, "prestige|NOUN": 4.9, "tolk|NOUN": 4.9, "reträtt|NOUN": 4.89, "nolla|NOUN": 4.89, "bricka|NOUN": 4.89, "korrigering|NOUN": 4.89, "lyxig|ADJ": 4.88, "reaktor|NOUN": 4.88, "banan|NOUN": 4.88, "kult|NOUN": 4.88, "komedi|NOUN": 4.87, "trick|NOUN": 4.87, "separation|NOUN": 4.86, "avlösa|VERB": 4.86, "betvivla|VERB": 4.86, "likaledes|ADV": 4.84, "retur|NOUN": 4.84, "dussin|NOUN": 4.84, "kylig|ADJ": 4.84, "dröjsmål|NOUN": 4.83, "grädde|NOUN": 4.83, "intellekt|NOUN": 4.83, "aggression|NOUN": 4.83, "buske|NOUN": 4.83, "minderårig|ADJ": 4.83, "spinna|VERB": 4.83, "interaktion|NOUN": 4.82, "terminologi|NOUN": 4.82, "östlig|ADJ": 4.82, "avsked|NOUN": 4.82, "hal|ADJ": 4.82, "rival|NOUN": 4.82, "proklamera|VERB": 4.81, "sofistikerad|ADJ": 4.81, "spruta|NOUN": 4.81, "anständig|ADJ": 4.8, "pump|NOUN": 4.8, "sexig|ADJ": 4.79, "förflyttning|NOUN": 4.78, "huvudsak|NOUN": 4.77, "utelämna|VERB": 4.77, "boskap|NOUN": 4.76, "exponera|VERB": 4.76, "lila|ADJ": 4.76, "tillägna|VERB": 4.76, "genus|NOUN": 4.76, "verb|NOUN": 4.76, "köpman|NOUN": 4.75, "vidarebefordra|VERB": 4.75, "frånta|VERB": 4.75, "interaktiv|ADJ": 4.75, "lagstifta|VERB": 4.75, "specialitet|NOUN": 4.75, "stråla|VERB": 4.75, "domkyrka|NOUN": 4.74, "slapp|ADJ": 4.74, "utvinna|VERB": 4.74, "upphöjd|ADJ": 4.73, "vykort|NOUN": 4.73, "assistans|NOUN": 4.73, "begåvning|NOUN": 4.73, "måleri|NOUN": 4.72, "påhitt|NOUN": 4.72, "kompakt|ADJ": 4.71, "samtycka|VERB": 4.71, "hälsovård|NOUN": 4.7, "lyft|NOUN": 4.7, "asfalt|NOUN": 4.7, "underkänna|VERB": 4.7, "uppoffring|NOUN": 4.7, "utrusta|VERB": 4.7, "förflyta|VERB": 4.69, "handledning|NOUN": 4.69, "oenighet|NOUN": 4.68, "slogan|NOUN": 4.68, "triumf|NOUN": 4.68, "färdigställa|VERB": 4.68, "skötsel|NOUN": 4.68, "portal|NOUN": 4.66, "överdrivet|ADV": 4.66, "applådera|VERB": 4.65, "husvagn|NOUN": 4.65, "vodka|NOUN": 4.65, "lansering|NOUN": 4.63, "handduk|NOUN": 4.63, "honung|NOUN": 4.62, "kanin|NOUN": 4.62, "målare|NOUN": 4.62, "plågsam|ADJ": 4.62, "trollkarl|NOUN": 4.61, "avancera|VERB": 4.61, "homogen|ADJ": 4.61, "skingra|VERB": 4.61, "underordna|VERB": 4.61, "överlägsenhet|NOUN": 4.61, "krocka|VERB": 4.6, "filt|NOUN": 4.59, "herravälde|NOUN": 4.59, "ryttare|NOUN": 4.59, "peppar|NOUN": 4.58, "nominell|ADJ": 4.58, "spola|VERB": 4.58, "defensiv|ADJ": 4.57, "katedral|NOUN": 4.57, "fjärran|ADJ": 4.56, "skär|ADJ": 4.56, "desperation|NOUN": 4.56, "blöda|VERB": 4.54, "ört|NOUN": 4.54, "avslappnad|ADJ": 4.54, "efterlevnad|NOUN": 4.53, "resande|NOUN": 4.53, "bär|NOUN": 4.51, "mysterium|NOUN": 4.51, "omvänt|ADV": 4.51, "lillasyster|NOUN": 4.5, "massage|NOUN": 4.5, "märkbar|ADJ": 4.49, "hane|NOUN": 4.49, "regelrätt|ADJ": 4.49, "gryning|NOUN": 4.48, "gudom|NOUN": 4.48, "överste|NOUN": 4.48, "uttråkad|ADJ": 4.48, "helikopter|NOUN": 4.47, "parasit|NOUN": 4.47, "utgrävning|NOUN": 4.47, "drake|NOUN": 4.47, "kryssa|VERB": 4.47, "stolpe|NOUN": 4.47, "kartong|NOUN": 4.46, "realism|NOUN": 4.46, "stackare|NOUN": 4.46, "höft|NOUN": 4.45, "skinka|NOUN": 4.45, "stökig|ADJ": 4.45, "råna|VERB": 4.45, "anförtro|VERB": 4.44, "försäljare|NOUN": 4.44, "gränssnitt|NOUN": 4.44, "stängning|NOUN": 4.44, "elfte|NUM": 4.43, "schack|NOUN": 4.43, "benägenhet|NOUN": 4.43, "intag|NOUN": 4.43, "stadion|NOUN": 4.42, "autentisk|ADJ": 4.41, "blankett|NOUN": 4.41, "fotografering|NOUN": 4.41, "rullstol|NOUN": 4.41, "årtal|NOUN": 4.41, "språng|NOUN": 4.4, "brunn|NOUN": 4.4, "artificiell|ADJ": 4.4, "företagsamhet|NOUN": 4.4, "filtrera|VERB": 4.39, "förolämpning|NOUN": 4.39, "kompani|NOUN": 0.6, "subventionera|VERB": 4.39, "uthållighet|NOUN": 4.39, "matsal|NOUN": 4.39, "skymning|NOUN": 4.38, "bekvämlighet|NOUN": 4.37, "eländig|ADJ": 4.37, "ark|NOUN": 3.3, "bulle|NOUN": 4.36, "parad|NOUN": 4.36, "stressa|VERB": 4.36, "glimt|NOUN": 4.36, "massaker|NOUN": 4.36, "riklig|ADJ": 4.35, "utlopp|NOUN": 4.35, "diplomati|NOUN": 4.34, "sås|NOUN": 4.34, "omfamna|VERB": 4.34, "absorbera|VERB": 4.33, "brandman|NOUN": 4.33, "lätthet|NOUN": 4.33, "uppslutning|NOUN": 4.33, "farväl|NOUN": 4.32, "specificera|VERB": 4.32, "broms|NOUN": 4.32, "dynasti|NOUN": 4.32, "tomrum|NOUN": 4.32, "förbrukning|NOUN": 4.32, "klia|VERB": 4.32, "tillgripa|VERB": 4.32, "trög|ADJ": 4.32, "välgörenhet|NOUN": 4.32, "instinkt|NOUN": 4.31, "hädanefter|ADV": 4.3, "utdela|VERB": 4.3, "adoption|NOUN": 4.3, "försvinnande|NOUN": 4.29, "gisslan|NOUN": 4.29, "kvalificera|VERB": 4.29, "nykomling|NOUN": 4.29, "prenumeration|NOUN": 4.28, "barack|NOUN": 4.28, "fotbollsspelare|NOUN": 4.28, "förevändning|NOUN": 4.28, "aha|INTJ": 4.27, "bukt|NOUN": 4.27, "grundtanke|NOUN": 4.27, "slicka|VERB": 4.27, "genial|ADJ": 4.26, "grind|NOUN": 4.26, "kuvert|NOUN": 4.26, "odödlig|ADJ": 4.26, "elektronik|NOUN": 4.26, "publicitet|NOUN": 4.25, "barnmorska|NOUN": 4.25, "påfallande|ADJ": 4.25, "kavaj|NOUN": 4.25, "lins|NOUN": 4.24, "psyke|NOUN": 4.23, "allergi|NOUN": 4.23, "resande|ADJ": 4.23, "specialisera|VERB": 4.23, "mognad|NOUN": 4.22, "skelett|NOUN": 4.22, "mager|ADJ": 4.21, "beslutsamhet|NOUN": 4.2, "brödraskap|NOUN": 4.19, "slumpmässig|ADJ": 4.19, "helgdag|NOUN": 4.18, "inlärning|NOUN": 4.18, "manuskript|NOUN": 4.18, "massvis|ADV": 4.18, "uppvisning|NOUN": 4.18, "följeslagare|NOUN": 4.18, "ovetande|ADJ": 4.18, "portfölj|NOUN": 4.18, "trohet|NOUN": 4.18, "kontant|ADJ": 4.18, "kontanter|NOUN": 4.18, "bomull|NOUN": 4.17, "höna|NOUN": 4.16, "nattvard|NOUN": 4.16, "rutt|NOUN": 4.16, "avsättning|NOUN": 4.15, "lår|NOUN": 4.15, "motbevisa|VERB": 4.15, "gröt|NOUN": 4.15, "logotyp|NOUN": 4.15, "nyårsafton|NOUN": 4.15, "fläkt|NOUN": 4.14, "högtalare|NOUN": 4.14, "kräkas|VERB": 4.13, "lokalisera|VERB": 4.13, "lantbruk|NOUN": 4.13, "fjäril|NOUN": 4.11, "officer|NOUN": 4.11, "påbud|NOUN": 4.11, "underkläder|NOUN": 4.11, "hastig|ADJ": 4.11, "faster|NOUN": 4.11, "sammankalla|VERB": 4.11, "anekdot|NOUN": 4.11, "rekommenderad|ADJ": 4.11, "dike|NOUN": 4.1, "parfym|NOUN": 4.1, "intuition|NOUN": 4.08, "kortvarig|ADJ": 4.08, "växthus|NOUN": 4.08, "modul|NOUN": 4.07, "fantisera|VERB": 4.06, "landsman|NOUN": 4.06, "skönlitteratur|NOUN": 4.06, "maka|NOUN": 4.06, "prosa|NOUN": 4.05, "användbarhet|NOUN": 4.05, "förläggare|NOUN": 4.05, "förolämpa|VERB": 4.05, "påföljande|ADJ": 4.05, "notering|NOUN": 4.04, "nål|NOUN": 4.04, "talrik|ADJ": 4.04, "komplettering|NOUN": 4.03, "ordspråk|NOUN": 4.03, "solnedgång|NOUN": 4.03, "attribut|NOUN": 4.01, "fosterland|NOUN": 4.01, "klot|NOUN": 4.01, "utbetala|VERB": 4.01, "alfabet|NOUN": 3.99, "bokföring|NOUN": 3.99, "fräck|ADJ": 3.99, "gammaldags|ADJ": 3.99, "Jorden|PROPN": 3.99, "jaså|INTJ": 3.98, "lämplighet|NOUN": 3.98, "sönderfall|NOUN": 3.98, "ämbetsman|NOUN": 3.98, "duell|NOUN": 3.97, "likviditet|NOUN": 3.97, "lossna|VERB": 3.97, "mikrofon|NOUN": 3.97, "trottoar|NOUN": 3.97, "slips|NOUN": 3.97, "hormon|NOUN": 3.96, "illamående|NOUN": 3.96, "tilldelning|NOUN": 3.96, "aluminium|NOUN": 3.96, "kappa|NOUN": 3.96, "permission|NOUN": 3.96, "försprång|NOUN": 3.95, "intim|ADJ": 3.95, "älskare|NOUN": 3.95, "skvaller|NOUN": 3.95, "metodik|NOUN": 3.94, "attraktion|NOUN": 3.94, "fragment|NOUN": 3.94, "magister|NOUN": 3.94, "reserv|NOUN": 3.94, "ekologi|NOUN": 3.93, "sponsring|NOUN": 3.92, "adelsman|NOUN": 3.91, "maskineri|NOUN": 3.91, "spalt|NOUN": 3.91, "underkastelse|NOUN": 3.9, "uråldrig|ADJ": 3.9, "clown|NOUN": 3.9, "noll|NOUN": 3.9, "verbal|ADJ": 3.9, "framträdande|NOUN": 3.89, "polisstation|NOUN": 3.89, "borsta|VERB": 3.89, "bägare|NOUN": 3.89, "gränslös|ADJ": 3.89, "kärl|NOUN": 3.88, "utomordentlig|ADJ": 3.88, "manager|NOUN": 3.88, "sångerska|NOUN": 3.88, "kooperativ|NOUN": 3.87, "genomskinlig|ADJ": 3.86, "kalender|NOUN": 3.85, "option|NOUN": 3.85, "arkeolog|NOUN": 3.85, "oändlighet|NOUN": 3.84, "netto|NOUN": 3.84, "veto|NOUN": 3.84, "veteran|NOUN": 3.82, "kalori|NOUN": 3.81, "vits|NOUN": 3.81, "kruka|NOUN": 3.8, "lotteri|NOUN": 3.8, "spektrum|NOUN": 3.8, "attentat|NOUN": 3.8, "avtala|VERB": 3.8, "förutsägelse|NOUN": 3.79, "halvtid|NOUN": 3.79, "kvitto|NOUN": 3.78, "oförutsedd|ADJ": 3.77, "livskraftig|ADJ": 3.77, "delegera|VERB": 3.76, "flit|NOUN": 3.76, "fullvärdig|ADJ": 3.75, "stab|NOUN": 3.75, "päron|NOUN": 3.75, "myndig|ADJ": 3.75, "förräderi|NOUN": 3.74, "förskott|NOUN": 3.74, "raka|VERB": 3.74, "svida|VERB": 3.74, "syntetisk|ADJ": 3.74, "mala|VERB": 3.73, "frisör|NOUN": 3.73, "osanning|NOUN": 3.73, "identifiering|NOUN": 3.72, "undre|ADJ": 3.72, "återvinning|NOUN": 3.72, "hurra|VERB": 3.71, "landning|NOUN": 3.71, "spilla|VERB": 3.71, "duva|NOUN": 3.71, "pryda|VERB": 3.71, "karakterisera|VERB": 3.7, "komponera|VERB": 3.7, "vidsträckt|ADJ": 3.7, "areal|NOUN": 3.69, "utvecklare|NOUN": 3.69, "betjäna|VERB": 3.69, "projektion|NOUN": 3.69, "skrattretande|ADJ": 3.69, "bacon|NOUN": 3.68, "gräl|NOUN": 3.68, "diameter|NOUN": 3.68, "förhöra|VERB": 3.68, "läsk|NOUN": 3.68, "tillmäta|VERB": 3.68, "åsna|NOUN": 3.67, "konsolidering|NOUN": 3.67, "tidtabell|NOUN": 3.67, "återbetalning|NOUN": 3.67, "explicit|ADV": 3.66, "kafé (el. café)|NOUN": 3.66, "manifest|ADJ": 3.66, "stram|ADJ": 3.66, "handske|NOUN": 3.65, "informativ|ADJ": 3.65, "rekonstruktion|NOUN": 3.65, "ridning|NOUN": 3.65, "garn|NOUN": 3.65, "samtidig|ADJ": 3.64, "matt|ADJ": 3.64, "bredda|VERB": 3.63, "gruppledare|NOUN": 3.63, "certifikat|NOUN": 3.62, "garage|NOUN": 3.62, "sociologi|NOUN": 3.62, "angränsande|ADJ": 3.61, "festlig|ADJ": 3.61, "generalisera|VERB": 3.61, "glödlampa|NOUN": 3.61, "grubbla|VERB": 3.61, "lantbrukare|NOUN": 3.61, "stipendium|NOUN": 3.61, "strukturera|VERB": 3.61, "tjur|NOUN": 3.61, "böna|NOUN": 3.61, "erotisk|ADJ": 3.6, "förträfflig|ADJ": 3.59, "löpare|NOUN": 3.59, "medlidande|NOUN": 3.59, "spänd|ADJ": 3.58, "gardin|NOUN": 3.58, "programmerare|NOUN": 3.58, "radiostation|NOUN": 3.58, "hosta|VERB": 3.57, "jämvikt|NOUN": 3.57, "tonvikt|NOUN": 3.57, "lobby|NOUN": 3.57, "explosiv|ADJ": 3.56, "hjälplös|ADJ": 3.56, "klausul|NOUN": 3.56, "spindel|NOUN": 3.55, "topplista|NOUN": 3.55, "klump|NOUN": 3.55, "trivsam|ADJ": 3.54, "brådskande|ADJ": 3.54, "elementär|ADJ": 3.54, "rättfärdiga|VERB": 3.54, "navigera|VERB": 3.54, "darra|VERB": 3.53, "flygel|NOUN": 3.53, "orientering|NOUN": 3.53, "utpräglad|ADJ": 3.53, "bebo|VERB": 3.53, "embryo|NOUN": 3.53, "lexikon|NOUN": 3.53, "experimentell|ADJ": 3.52, "instifta|VERB": 3.52, "väsentligen|ADV": 3.52, "kortfattad|ADJ": 3.52, "referat|NOUN": 3.52, "fyr|NOUN": 3.51, "förbränning|NOUN": 3.51, "inrymma|VERB": 3.51, "privilegierad|ADJ": 3.51, "kardinal|NOUN": 3.5, "essens|NOUN": 3.5, "affärsverksamhet|NOUN": 3.48, "extraordinär|ADJ": 3.48, "grammatik|NOUN": 3.48, "komposition|NOUN": 3.48, "krok|NOUN": 3.48, "kyss|NOUN": 3.47, "företrädesvis|ADV": 3.47, "medfödd|ADJ": 3.47, "jurisdiktion|NOUN": 3.46, "knipa|VERB": 3.46, "kondition|NOUN": 3.46, "oriktig|ADJ": 3.46, "proportionell|ADJ": 3.46, "själslig|ADJ": 3.46, "dagsljus|NOUN": 3.46, "fukt|NOUN": 3.46, "abonnemang|NOUN": 3.45, "sammanföra|VERB": 3.45, "ånga|NOUN": 3.45, "aktiemarknad|NOUN": 3.44, "mapp|NOUN": 3.44, "prototyp|NOUN": 3.44, "vilseleda|VERB": 3.44, "immigrant|NOUN": 3.43, "anlag|NOUN": 3.43, "fullmakt|NOUN": 3.43, "hyresvärd|NOUN": 3.43, "klassificering|NOUN": 3.43, "parlamentsledamot|NOUN": 3.43, "försena|VERB": 3.42, "renhet|NOUN": 3.41, "övertid|NOUN": 3.41, "allergisk|ADJ": 3.4, "eskalera|VERB": 3.4, "föreståndare|NOUN": 3.4, "spanare|NOUN": 3.4, "instruktör|NOUN": 3.4, "mugg|NOUN": 3.4, "granat|NOUN": 3.4, "ofrivillig|ADJ": 3.39, "subtil|ADJ": 3.39, "successiv|ADJ": 3.39, "välvilja|NOUN": 3.39, "banal|ADJ": 3.39, "spjut|NOUN": 3.39, "hektar|NOUN": 3.39, "avvärja|VERB": 3.38, "hållplats|NOUN": 3.38, "härma|VERB": 3.38, "distributör|NOUN": 3.37, "hårdvara|NOUN": 3.36, "grop|NOUN": 3.36, "repetera|VERB": 3.36, "utrotning|NOUN": 3.36, "grannskap|NOUN": 3.35, "kamel|NOUN": 3.35, "avlopp|NOUN": 3.35, "hjälpsam|ADJ": 3.35, "ämnesområde|NOUN": 3.35, "ändlös|ADJ": 3.35, "flamma|NOUN": 3.35, "livmoder|NOUN": 3.34, "reduktion|NOUN": 3.34, "susa|VERB": 3.34, "funktionalitet|NOUN": 3.33, "kulminera|VERB": 3.33, "slät|ADJ": 3.33, "hysteri|NOUN": 3.33, "rulle|NOUN": 3.33, "nattlig|ADJ": 3.32, "stråle|NOUN": 3.32, "avskilja|VERB": 3.32, "värdesätta|VERB": 3.32, "bark|NOUN": 3.31, "nalle|NOUN": 3.31, "fångst|NOUN": 3.31, "revolutionerande|ADJ": 3.31, "fåtölj|NOUN": 3.3, "ogiltig|ADJ": 3.3, "hygien|NOUN": 3.3, "tegel|NOUN": 3.3, "accelerera|VERB": 3.29, "gedigen|ADJ": 3.28, "känslighet|NOUN": 3.28, "sluttning|NOUN": 3.28, "nordväst|NOUN": 3.27, "utsökt|ADJ": 3.27, "analogi|NOUN": 3.27, "specifikation|NOUN": 3.27, "samordnare|NOUN": 3.26, "stöt|NOUN": 3.26, "bandit|NOUN": 3.26, "devalvering|NOUN": 3.25, "internationalisering|NOUN": 3.25, "kölvatten|NOUN": 3.25, "frige|VERB": 3.25, "åska|NOUN": 3.25, "hallå|NOUN": 3.25, "badkar|NOUN": 3.25, "obligation|NOUN": 3.25, "vertikal|ADJ": 3.25, "sommarlov|NOUN": 3.23, "volontär|NOUN": 3.23, "likgiltighet|NOUN": 3.23, "mottaglig|ADJ": 3.23, "noggrannhet|NOUN": 3.23, "tjat|NOUN": 3.23, "addera|VERB": 3.21, "barnvagn|NOUN": 3.21, "hurra|INTJ": 3.21, "simning|NOUN": 3.21, "omvårdnad|NOUN": 3.21, "beskydda|VERB": 3.2, "fyrkantig|ADJ": 3.2, "tunna|NOUN": 3.2, "ull|NOUN": 3.2, "avresa|NOUN": 3.19, "båge|NOUN": 3.19, "robust|ADJ": 3.19, "suppleant|NOUN": 3.19, "energisk|ADJ": 3.19, "rikligt|ADV": 3.19, "blotta|VERB": 3.18, "lokalisering|NOUN": 3.18, "interagera|VERB": 3.18, "julgran|NOUN": 3.18, "porto|NOUN": 3.18, "stick|NOUN": 3.17, "rotera|VERB": 3.17, "kiosk|NOUN": 3.16, "galler|NOUN": 3.16, "onormal|ADJ": 3.15, "oräknelig|ADJ": 3.15, "olivolja|NOUN": 3.15, "bokning|NOUN": 3.14, "förskräcklig|ADJ": 3.14, "inspektera|VERB": 3.14, "orientera|VERB": 3.14, "smeka|VERB": 3.14, "välgörande|ADJ": 3.14, "reception|NOUN": 3.14, "reproduktion|NOUN": 3.13, "konsul|NOUN": 3.12, "konsulat|NOUN": 3.12, "medvetslös|ADJ": 3.12, "moped|NOUN": 3.12, "sammanträda|VERB": 3.12, "altare|NOUN": 3.11, "kidnappning|NOUN": 3.11, "uppfyllelse|NOUN": 3.11, "betingelse|NOUN": 3.11, "förplikta|VERB": 3.11, "handväska|NOUN": 3.11, "häkta|VERB": 3.11, "rådjur|NOUN": 3.11, "specialisering|NOUN": 3.11, "överfall|NOUN": 3.11, "frimärke|NOUN": 3.1, "lakan|NOUN": 3.1, "gurka|NOUN": 3.09, "kanna|NOUN": 3.09, "midja|NOUN": 3.09, "omringa|VERB": 3.09, "styrelseordförande|NOUN": 3.09, "ödelägga|VERB": 3.09, "slang|NOUN": 3.08, "överhuvud|NOUN": 3.08, "handelsman|NOUN": 3.08, "linjär|ADJ": 3.08, "telekommunikation|NOUN": 3.08, "karakteristisk|ADJ": 3.07, "åklagarmyndighet|NOUN": 3.07, "årsdag|NOUN": 3.07, "repetition|NOUN": 3.07, "underskrift|NOUN": 3.06, "förgrund|NOUN": 3.05, "grönska|NOUN": 3.05, "kungörelse|NOUN": 3.05, "besvära|VERB": 3.04, "reflex|NOUN": 3.04, "inspektör|NOUN": 3.04, "stum|ADJ": 3.04, "uppdra|VERB": 3.04, "gunga|VERB": 3.04, "kooperativ|ADJ": 3.04, "legitimation|NOUN": 3.04, "patriotisk|ADJ": 3.04, "aptit|NOUN": 3.03, "artig|ADJ": 3.03, "beskyddare|NOUN": 3.03, "samstämmighet|NOUN": 3.03, "uppehälle|NOUN": 3.03, "segment|NOUN": 3.03, "stege|NOUN": 3.03, "rea|NOUN": 3.02, "oliv|NOUN": 3.01, "syra|NOUN": 3.01, "vattna|VERB": 3.01, "besätta|VERB": 3.01, "dispyt|NOUN": 3.01, "kräfta|NOUN": 3.0, "läcker|ADJ": 3.0, "vaktmästare|NOUN": 3.0, "byggnation|NOUN": 2.99, "förlåt|INTJ": 2.99, "bi|NOUN": 2.99, "dårskap|NOUN": 2.99, "räka|NOUN": 2.99, "terminal|NOUN": 2.98, "vakuum|NOUN": 2.98, "fusion|NOUN": 2.97, "utskrift|NOUN": 2.97, "offert|NOUN": 2.97, "botemedel|NOUN": 2.96, "säregen|ADJ": 2.96, "taxa|NOUN": 2.96, "välvillig|ADJ": 2.96, "klumpig|ADJ": 2.96, "tillflykt|NOUN": 2.96, "vävnad|NOUN": 2.96, "majestät|NOUN": 2.96, "immunitet|NOUN": 2.95, "ombildning|NOUN": 2.95, "omstridd|ADJ": 2.95, "periferi|NOUN": 2.95, "nunna|NOUN": 2.95, "löjtnant|NOUN": 2.94, "återlämna|VERB": 2.94, "stav|NOUN": 2.93, "fridfull|ADJ": 2.93, "höghus|NOUN": 2.93, "innevånare|NOUN": 2.93, "sjösätta|VERB": 2.93, "trauma|NOUN": 2.93, "oväder|NOUN": 2.92, "spion|NOUN": 2.92, "komplicera|VERB": 2.92, "substantiv|NOUN": 2.92, "undersida|NOUN": 2.92, "putsa|VERB": 2.91, "kam|NOUN": 2.91, "manuell|ADJ": 2.91, "mittfält|NOUN": 2.91, "pizzeria|NOUN": 2.91, "sittplats|NOUN": 2.9, "uthyrning|NOUN": 2.9, "komplimang|NOUN": 2.9, "handtag|NOUN": 2.9, "bemästra|VERB": 2.89, "obekant|ADJ": 2.89, "stapla|VERB": 2.89, "tusental|NOUN": 2.89, "berättiga|VERB": 2.89, "stereotyp|ADJ": 2.89, "vitlök|NOUN": 2.88, "alkoholism|NOUN": 2.87, "beröring|NOUN": 2.87, "bete|NOUN": 2.87, "flerårig|ADJ": 2.87, "förråda|VERB": 2.87, "försändelse|NOUN": 2.87, "resväska|NOUN": 2.87, "flyktig|ADJ": 2.86, "kirurg|NOUN": 2.86, "otvivelaktigt|ADV": 2.86, "saft|NOUN": 2.86, "varaktighet|NOUN": 2.86, "lekplats|NOUN": 2.85, "tillförlitlighet|NOUN": 2.85, "adjö|INTJ": 2.84, "käpp|NOUN": 2.84, "lossa|VERB": 2.84, "summering|NOUN": 2.84, "exekutiv|ADJ": 2.83, "kandidatur|NOUN": 2.83, "tum|NOUN": 2.83, "återkoppling|NOUN": 2.83, "dofta|VERB": 2.82, "encyklopedi|NOUN": 2.82, "förrädare|NOUN": 2.82, "tvättmaskin|NOUN": 2.82, "kvist|NOUN": 2.82, "tvål|NOUN": 2.82, "madrass|NOUN": 2.82, "heder|NOUN": 2.81, "knop|NOUN": 2.81, "maträtt|NOUN": 2.81, "njure|NOUN": 2.81, "alstra|VERB": 2.81, "beslutsam|ADJ": 2.81, "kontur|NOUN": 2.81, "värka|VERB": 2.81, "droppe|NOUN": 2.8, "inställa|VERB": 2.8, "programmera|VERB": 2.8, "resebyrå|NOUN": 2.8, "gnista|NOUN": 2.8, "envishet|NOUN": 2.79, "stilig|ADJ": 2.79, "vänskaplig|ADJ": 2.79, "kristall|NOUN": 2.78, "passionerad|ADJ": 2.78, "yr|ADJ": 2.78, "besiktning|NOUN": 2.78, "delgivning|NOUN": 2.78, "gjuta|VERB": 2.78, "smörja|VERB": 2.78, "ådra|VERB": 2.78, "åkomma|NOUN": 2.78, "stång|NOUN": 2.77, "konsultera|VERB": 2.77, "återuppliva|VERB": 2.77, "växtlighet|NOUN": 2.76, "frost|NOUN": 2.76, "lykta|NOUN": 2.76, "akustisk|ADJ": 2.75, "antydning|NOUN": 2.75, "häl|NOUN": 2.75, "hängivenhet|NOUN": 2.75, "orätt|NOUN": 2.75, "syntes|NOUN": 2.75, "ungdomlig|ADJ": 2.75, "citron|NOUN": 2.75, "tillbakadragande|NOUN": 2.75, "förfalskning|NOUN": 2.75, "tass|NOUN": 2.75, "trasa|NOUN": 2.75, "orgel|NOUN": 2.74, "oberoende|NOUN": 2.74, "geometri|NOUN": 2.73, "omfång|NOUN": 2.73, "oviss|ADJ": 2.73, "uteslutning|NOUN": 2.73, "utsända|VERB": 2.73, "pensionering|NOUN": 2.72, "förstora|VERB": 2.72, "försvinnande|ADV": 2.72, "paraply|NOUN": 2.72, "plakat|NOUN": 2.72, "veranda|NOUN": 2.72, "kosttillskott|NOUN": 2.71, "krock|NOUN": 2.71, "skyltfönster|NOUN": 2.71, "munter|ADJ": 2.71, "shorts|NOUN": 2.71, "vandrarhem|NOUN": 2.71, "kvadrat|NOUN": 2.7, "raseri|NOUN": 2.7, "tangent|NOUN": 2.7, "interiör|NOUN": 2.69, "bondgård|NOUN": 2.69, "brådska|NOUN": 2.69, "svartsjuka|NOUN": 2.69, "älskarinna|NOUN": 2.69, "adjektiv|NOUN": 2.68, "berömmelse|NOUN": 2.68, "bundsförvant|NOUN": 2.68, "fjärran|ADV": 2.68, "utantill|ADV": 2.68, "överträda|VERB": 2.68, "bortskämd|ADJ": 2.68, "byggare|NOUN": 2.68, "obildad|ADJ": 2.68, "bål|NOUN": 0.68, "horisontell|ADJ": 2.68, "imitera|VERB": 2.68, "optisk|ADJ": 2.68, "temperament|NOUN": 2.68, "uppställning|NOUN": 2.68, "bedragare|NOUN": 2.67, "tonfall|NOUN": 2.67, "fotografisk|ADJ": 2.66, "skissera|VERB": 2.66, "kollision|NOUN": 2.65, "magnetisk|ADJ": 2.64, "sparsam|ADJ": 2.64, "prestigefylld|ADJ": 2.64, "kran|NOUN": 2.63, "småstad|NOUN": 2.63, "vingård|NOUN": 2.63, "flamma|VERB": 2.62, "försona|VERB": 2.62, "treårig|ADJ": 2.62, "utlämna|VERB": 2.62, "linne|NOUN": 2.61, "nybyggare|NOUN": 2.61, "triangel|NOUN": 2.61, "utsliten|ADJ": 2.61, "slank|ADJ": 2.61, "annullera|VERB": 2.6, "brandkår|NOUN": 2.6, "pinne|NOUN": 2.6, "hare|NOUN": 2.6, "jämförande|ADJ": 2.6, "ministerium|NOUN": 2.6, "vikarie|NOUN": 2.59, "astma|NOUN": 2.59, "förvirra|VERB": 2.59, "inflammation|NOUN": 2.59, "larma|VERB": 2.59, "mätta|VERB": 2.59, "plåster|NOUN": 2.58, "rotation|NOUN": 2.58, "skolgård|NOUN": 2.58, "åtkomst|NOUN": 2.58, "övernatta|VERB": 2.58, "egenhet|NOUN": 2.57, "oordning|NOUN": 2.57, "revidering|NOUN": 2.57, "smörja|NOUN": 2.57, "ålderdom|NOUN": 2.57, "kommando|NOUN": 2.57, "utmattning|NOUN": 2.56, "keramik|NOUN": 2.56, "mustasch|NOUN": 2.56, "baron|NOUN": 2.55, "boss|NOUN": 2.55, "läder|NOUN": 2.55, "rengöring|NOUN": 2.55, "avfärd|NOUN": 2.55, "hink|NOUN": 2.55, "matematiker|NOUN": 2.55, "passning|NOUN": 2.55, "tillsättning|NOUN": 2.55, "hemort|NOUN": 2.54, "instruera|VERB": 2.54, "rengöra|VERB": 2.54, "dekoration|NOUN": 2.54, "månatlig|ADJ": 2.54, "patriotism|NOUN": 2.54, "tillmötesgå|VERB": 2.54, "gås|NOUN": 2.54, "programmering|NOUN": 2.53, "vicepresident|NOUN": 2.53, "avla|VERB": 2.53, "brigad|NOUN": 2.53, "allsidig|ADJ": 2.52, "komfort|NOUN": 2.52, "listig|ADJ": 2.52, "simulering|NOUN": 2.52, "återbetala|VERB": 2.52, "sned|ADJ": 2.51, "bassäng|NOUN": 2.51, "närbelägen|ADJ": 2.51, "pensel|NOUN": 2.51, "luftfart|NOUN": 2.5, "patrull|NOUN": 2.5, "arbetsrum|NOUN": 2.5, "implementering|NOUN": 2.5, "hydda|NOUN": 2.49, "oerfaren|ADJ": 2.49, "bokstavlig|ADJ": 2.47, "elektromagnetisk|ADJ": 2.47, "rymlig|ADJ": 2.47, "världsåskådning|NOUN": 2.46, "ansiktsuttryck|NOUN": 2.46, "frigivning|NOUN": 2.46, "pristagare|NOUN": 2.46, "självsäker|ADJ": 2.46, "fiber|NOUN": 2.46, "dricks|NOUN": 2.45, "tam|ADJ": 2.45, "oreda|NOUN": 2.44, "förnekande|NOUN": 2.43, "algoritm|NOUN": 2.42, "tall|NOUN": 2.42, "avsiktlig|ADJ": 2.42, "biolog|NOUN": 2.42, "tarm|NOUN": 2.42, "adlig|ADJ": 2.41, "spegelbild|NOUN": 2.41, "campus|NOUN": 2.41, "brännvin|NOUN": 2.4, "kompatibel|ADJ": 2.4, "ängslig|ADJ": 2.4, "tolfte|NUM": 2.4, "beväpna|VERB": 2.4, "tvåhundra|NUM": 2.4, "biff|NOUN": 2.39, "ratificering|NOUN": 2.39, "skådespelerska|NOUN": 2.39, "slavisk|ADJ": 2.39, "glänsa|VERB": 2.39, "ömhet|NOUN": 2.39, "föräldralös|ADJ": 2.38, "tumör|NOUN": 2.38, "vidareutveckling|NOUN": 2.38, "juice|NOUN": 2.38, "deponera|VERB": 2.37, "kirurgi|NOUN": 2.37, "närmande|NOUN": 2.37, "rondell|NOUN": 2.37, "sensationell|ADJ": 2.37, "stabilisering|NOUN": 2.37, "törst|NOUN": 2.36, "arkitektonisk|ADJ": 2.36, "förbluffande|ADV": 2.36, "klunga|NOUN": 2.36, "medfölja|VERB": 2.36, "processor|NOUN": 2.36, "tabu|ADJ": 2.36, "vulgär|ADJ": 2.36, "minnesmärke|NOUN": 2.35, "provision|NOUN": 2.35, "blödning|NOUN": 2.34, "defekt|NOUN": 2.34, "disposition|NOUN": 2.34, "koordinera|VERB": 2.34, "staket|NOUN": 2.34, "hytt|NOUN": 2.33, "kastrull|NOUN": 2.33, "startpunkt|NOUN": 2.33, "sked|NOUN": 2.33, "bal|NOUN": 2.33, "sandstrand|NOUN": 2.32, "stereotyp|NOUN": 2.32, "tålmodigt|ADV": 2.32, "arrestering|NOUN": 2.31, "kryssning|NOUN": 2.31, "pipa|VERB": 2.31, "gräla|VERB": 2.3, "area|NOUN": 2.3, "förbipasserande|ADJ": 2.3, "förlikning|NOUN": 2.29, "ljuda|VERB": 2.29, "samexistens|NOUN": 2.29, "terapeutisk|ADJ": 2.29, "trendig|ADJ": 2.29, "återhållsamhet|NOUN": 2.29, "hjort|NOUN": 2.29, "debitera|VERB": 2.28, "dundra|VERB": 2.28, "kräm|NOUN": 2.28, "korrespondent|NOUN": 2.27, "aktualitet|NOUN": 2.27, "behållare|NOUN": 2.26, "gruvarbetare|NOUN": 2.26, "åtstramning|NOUN": 2.26, "kontinental|ADJ": 2.26, "väster|NOUN": 2.26, "ankare|NOUN": 2.25, "åker|NOUN": 2.25, "senator|NOUN": 2.25, "häpnad|NOUN": 2.25, "mynning|NOUN": 2.25, "omtänksam|ADJ": 2.25, "omåttlig|ADJ": 2.25, "rekonstruera|VERB": 2.25, "maximum|NOUN": 2.24, "karaktärsdrag|NOUN": 2.23, "perfektion|NOUN": 2.23, "timmer|NOUN": 2.23, "urin|NOUN": 2.23, "arkivera|VERB": 2.22, "oavbruten|ADJ": 2.22, "kolonn|NOUN": 2.21, "appell|NOUN": 2.2, "strejka|VERB": 2.2, "propp|NOUN": 2.2, "automat|NOUN": 2.19, "studium|NOUN": 2.19, "högljudd|ADJ": 2.19, "skaldjur|NOUN": 2.19, "stinka|VERB": 2.19, "tillfreds|ADJ": 2.19, "världsomfattande|ADJ": 2.19, "befruktning|NOUN": 2.18, "glänsande|ADJ": 2.18, "organisatör|NOUN": 2.18, "pussel|NOUN": 2.18, "vitamin|NOUN": 2.18, "aktning|NOUN": 2.18, "boplats|NOUN": 2.18, "vederbörlig|ADJ": 2.18, "dråp|NOUN": 2.17, "jubileum|NOUN": 2.17, "frikänna|VERB": 2.17, "hetta|VERB": 2.17, "formation|NOUN": 2.16, "ridå|NOUN": 2.16, "rådfråga|VERB": 2.16, "svälla|VERB": 2.16, "avföring|NOUN": 2.15, "modifikation|NOUN": 2.14, "ordförråd|NOUN": 2.14, "tjocklek|NOUN": 2.14, "metropol|NOUN": 2.13, "injektion|NOUN": 2.13, "lantlig|ADJ": 2.13, "veckotidning|NOUN": 2.12, "orkester|NOUN": 2.11, "skruv|NOUN": 2.11, "solsken|NOUN": 2.11, "matvara|NOUN": 2.11, "regemente|NOUN": 2.11, "sammanträffande|NOUN": 2.11, "utstrålning|NOUN": 2.11, "valla|VERB": 2.11, "arvode|NOUN": 2.11, "periodisk|ADJ": 2.11, "favör|NOUN": 2.1, "kommunikativ|ADJ": 2.1, "terminal|ADJ": 2.1, "trappsteg|NOUN": 2.1, "paj|NOUN": 2.09, "anskaffa|VERB": 2.09, "mörkhyad|ADJ": 2.08, "tristess|NOUN": 2.08, "kassett|NOUN": 2.08, "räddare|NOUN": 2.08, "almanacka|NOUN": 2.07, "accent|NOUN": 2.07, "kvällsmat|NOUN": 2.07, "bestiga|VERB": 2.06, "styv|ADJ": 2.05, "knekt|NOUN": 2.05, "väv|NOUN": 2.05, "översvämma|VERB": 2.05, "örn|NOUN": 2.04, "seglare|NOUN": 2.04, "spöke|NOUN": 2.04, "lund|NOUN": 2.04, "tålmodig|ADJ": 2.04, "koja|NOUN": 2.03, "lockelse|NOUN": 2.03, "lärd|ADJ": 2.03, "balk|NOUN": 2.03, "åldring|NOUN": 2.02, "fullmåne|NOUN": 2.01, "bröstkorg|NOUN": 2.01, "slätt|ADV": 2.01, "spektakel|NOUN": 2.0, "ven|NOUN": 2.0, "nöt|NOUN": 2.0, "odjur|NOUN": 2.0, "äventyrare|NOUN": 2.0, "bildlig|ADJ": 1.99, "rangordna|VERB": 1.99, "smörgås|NOUN": 1.99, "hjord|NOUN": 1.99, "vildsvin|NOUN": 1.98, "bibliografi|NOUN": 1.97, "ihärdig|ADJ": 1.97, "indignation|NOUN": 1.97, "paradoxal|ADJ": 1.97, "soluppgång|NOUN": 1.97, "grädda|VERB": 1.97, "kontrovers|NOUN": 1.96, "multiplicera|VERB": 1.96, "oförrätt|NOUN": 1.96, "revben|NOUN": 1.96, "yoghurt|NOUN": 1.96, "delikat|ADJ": 1.95, "konsultation|NOUN": 1.95, "kväve|NOUN": 1.95, "kvarn|NOUN": 1.95, "gummi|NOUN": 1.94, "facilitet|NOUN": 1.94, "mittemot (el. mitt emot)|ADP": 1.94, "oenig|ADJ": 1.94, "oföränderlig|ADJ": 1.94, "restaurering|NOUN": 1.94, "snuskig|ADJ": 1.94, "tågstation|NOUN": 1.94, "herde|NOUN": 1.93, "kål|NOUN": 1.93, "tillförsel|NOUN": 1.93, "avskrivning|NOUN": 1.92, "bemanning|NOUN": 1.92, "pytteliten|ADJ": 1.92, "cirkulation|NOUN": 1.91, "termisk|ADJ": 1.91, "ömtålig|ADJ": 1.91, "koda|VERB": 1.91, "kämpe|NOUN": 1.91, "besatthet|NOUN": 1.9, "fjärrkontroll|NOUN": 1.9, "juvel|NOUN": 1.9, "ponny|NOUN": 1.9, "bemanna|VERB": 1.9, "måtta|NOUN": 1.9, "dekorera|VERB": 1.89, "gaffel|NOUN": 1.89, "pilgrim|NOUN": 1.89, "ackumulera|VERB": 1.89, "getto|NOUN": 1.89, "skorsten|NOUN": 1.89, "antenn|NOUN": 1.88, "montering|NOUN": 1.88, "synbar|ADJ": 1.88, "vrå|NOUN": 1.88, "assistera|VERB": 1.87, "defensiv|NOUN": 1.87, "videokamera|NOUN": 1.87, "bataljon|NOUN": 1.87, "intelligens|NOUN": 1.87, "diplom|NOUN": 1.86, "konfiguration|NOUN": 1.86, "efterfölja|VERB": 1.86, "exemplarisk|ADJ": 1.86, "konsistens|NOUN": 1.86, "stelna|VERB": 1.86, "amortering|NOUN": 1.85, "avskrift|NOUN": 1.85, "bläck|NOUN": 1.85, "restaurera|VERB": 1.85, "pulver|NOUN": 1.84, "remsa|NOUN": 1.84, "apelsin|NOUN": 1.84, "cement|NOUN": 1.84, "trailer|NOUN": 1.84, "ljum|ADJ": 1.83, "sammanstötning|NOUN": 1.83, "stormig|ADJ": 1.83, "pina|NOUN": 1.83, "skift|NOUN": 1.83, "stöna|VERB": 1.83, "uppsyn|NOUN": 1.82, "återse|VERB": 1.82, "elektron|NOUN": 1.82, "oanvändbar|ADJ": 1.82, "sömnig|ADJ": 1.82, "emission|NOUN": 1.81, "omloppsbana|NOUN": 1.81, "blixtsnabbt|ADV": 1.81, "brevväxling|NOUN": 1.81, "ventil|NOUN": 1.81, "fresta|VERB": 1.8, "pekfinger|NOUN": 1.8, "sigill|NOUN": 1.8, "armbåge|NOUN": 1.79, "ljusblå|ADJ": 1.79, "skaft|NOUN": 1.79, "paviljong|NOUN": 1.78, "segerrik|ADJ": 1.77, "skenbar|ADJ": 1.77, "svartsjuk|ADJ": 1.77, "mångfaldig|ADJ": 1.76, "omlopp|NOUN": 1.76, "kemist|NOUN": 1.76, "dykning|NOUN": 1.75, "orörlig|ADJ": 1.75, "tagning|NOUN": 1.75, "cykelväg|NOUN": 1.75, "donator|NOUN": 1.75, "förverkligande|NOUN": 1.75, "nyck|NOUN": 1.75, "gränsområde|NOUN": 1.74, "pittoresk|ADJ": 1.74, "yla|VERB": 1.74, "disciplinär|ADJ": 1.73, "farväl|INTJ": 1.73, "pånyttfödelse|NOUN": 1.73, "relik|NOUN": 1.73, "berättigande|NOUN": 1.72, "föresats|NOUN": 1.72, "inbetalning|NOUN": 1.72, "ströva|VERB": 1.72, "substitut|NOUN": 1.72, "tjugonde|NUM": 1.72, "arbetslag|NOUN": 1.72, "lim|NOUN": 1.72, "läglig|ADJ": 1.71, "nyttighet|NOUN": 1.71, "simhall|NOUN": 1.71, "animation|NOUN": 1.71, "väte|NOUN": 1.71, "orätt|ADJ": 1.7, "uppskov|NOUN": 1.7, "belägenhet|NOUN": 1.69, "sammandrag|NOUN": 1.69, "bensinstation|NOUN": 1.68, "gymnastik|NOUN": 1.68, "kommissarie|NOUN": 1.68, "vokal|NOUN": 1.68, "förmyndare|NOUN": 1.68, "mineral|NOUN": 1.68, "omnämnande|NOUN": 1.68, "alarm|NOUN": 1.67, "allé|NOUN": 1.67, "bergstopp|NOUN": 1.67, "navigation|NOUN": 1.67, "set|NOUN": 1.67, "tematisk|ADJ": 1.67, "täthet|NOUN": 1.67, "återupptäcka|VERB": 1.67, "postkontor|NOUN": 1.66, "ärm|NOUN": 1.65, "residens|NOUN": 1.65, "teleskop|NOUN": 1.65, "tryckning|NOUN": 1.64, "drickande|NOUN": 1.64, "kabinett|NOUN": 1.63, "charmerande|ADJ": 1.63, "missfall|NOUN": 1.63, "äktenskaplig|ADJ": 1.63, "emigrant|NOUN": 1.62, "bagatell|NOUN": 1.62, "bestämdhet|NOUN": 1.62, "aveny|NOUN": 1.61, "hosta|NOUN": 1.61, "andedräkt|NOUN": 1.61, "bottenvåning|NOUN": 1.61, "förtrolig|ADJ": 1.61, "avskedande|NOUN": 1.6, "femtonde|NUM": 1.6, "avbetalning|NOUN": 1.59, "fotgängare|NOUN": 1.59, "lärarinna|NOUN": 1.59, "terrass|NOUN": 1.59, "monter|NOUN": 1.58, "sylt|NOUN": 1.58, "kila|VERB": 1.57, "tuggummi|NOUN": 1.57, "bildskärm|NOUN": 1.56, "eliminering|NOUN": 1.56, "kalkylera|VERB": 1.56, "agentur|NOUN": 1.56, "mellanliggande|ADJ": 1.56, "trosa|NOUN": 1.56, "såg|NOUN": 1.55, "fysiologisk|ADJ": 1.55, "uppfödning|NOUN": 1.55, "betinga|VERB": 1.54, "farförälder|NOUN": 1.54, "råolja|NOUN": 1.54, "ficklampa|NOUN": 1.54, "hårig|ADJ": 1.54, "tvättmedel|NOUN": 1.54, "förorena|VERB": 1.54, "marskalk|NOUN": 1.54, "böjning|NOUN": 1.53, "narkoman|NOUN": 1.53, "upphetsning|NOUN": 1.53, "uppköp|NOUN": 1.53, "mentor|NOUN": 1.53, "fyrverkeri|NOUN": 1.52, "kollegium|NOUN": 1.52, "spade|NOUN": 1.52, "differentiering|NOUN": 1.52, "infektera|VERB": 1.52, "veck|NOUN": 1.52, "limma|VERB": 1.51, "oväsen|NOUN": 1.51, "innesluta|VERB": 1.51, "klädesplagg|NOUN": 1.51, "musiker|NOUN": 1.51, "smaklös|ADJ": 1.51, "stigning|NOUN": 1.51, "bravo|INTJ": 1.5, "hjärtlig|ADJ": 1.5, "explicit|ADJ": 1.49, "idrottsman|NOUN": 1.49, "koncession|NOUN": 1.49, "ofördelaktig|ADJ": 1.49, "ädel|ADJ": 1.49, "epos|NOUN": 1.49, "fasta|NOUN": 1.48, "geting|NOUN": 1.48, "hedervärd|ADJ": 1.48, "hjältinna|NOUN": 1.48, "knipa|NOUN": 1.48, "frågeformulär|NOUN": 1.47, "densitet|NOUN": 1.47, "eskortera|VERB": 1.47, "rankning|NOUN": 1.47, "servitör|NOUN": 1.47, "svägerska|NOUN": 1.47, "förbrylla|VERB": 1.46, "skattemässig|ADJ": 1.46, "tillgivenhet|NOUN": 1.46, "avkomling|NOUN": 1.45, "diagnostisera|VERB": 1.45, "rådman|NOUN": 1.45, "sammanfoga|VERB": 1.45, "ögonkast|NOUN": 1.45, "designer|NOUN": 1.45, "basilika|NOUN": 1.44, "lem|NOUN": 1.44, "adressera|VERB": 1.44, "bagare|NOUN": 1.44, "veckoslut|NOUN": 1.44, "centrera|VERB": 1.43, "fotfolk|NOUN": 1.43, "fästmö|NOUN": 1.43, "illvilja|NOUN": 1.43, "inskrivning|NOUN": 1.43, "omkrets|NOUN": 1.42, "självdeklaration|NOUN": 1.42, "trehundra|NUM": 1.42, "logo|NOUN": 1.41, "fyndighet|NOUN": 1.4, "gästfrihet|NOUN": 1.4, "konfirmation|NOUN": 1.4, "skär|NOUN": 1.4, "vindruva|NOUN": 1.4, "vårdare|NOUN": 1.4, "ådra|NOUN": 1.4, "tillfredsställd|ADJ": 1.4, "förestå|VERB": 1.39, "handflata|NOUN": 1.39, "inbillning|NOUN": 1.39, "logg|NOUN": 1.39, "bakverk|NOUN": 1.39, "gratulation|NOUN": 1.39, "kapplöpning|NOUN": 1.39, "opponent|NOUN": 1.39, "betydlig|ADJ": 1.38, "matris|NOUN": 1.38, "avdela|VERB": 1.37, "huvudämne|NOUN": 1.37, "komplott|NOUN": 1.37, "returnera|VERB": 1.37, "stadfästa|VERB": 1.37, "oavgjord|ADJ": 1.36, "beslutsamt|ADV": 1.36, "kupong|NOUN": 1.36, "massera|VERB": 1.36, "tändsticka|NOUN": 1.36, "ädelsten|NOUN": 1.36, "kakao|NOUN": 1.35, "akvarium|NOUN": 1.34, "smycke|NOUN": 1.34, "försvarsadvokat|NOUN": 1.33, "knytnäve|NOUN": 1.33, "optik|NOUN": 1.33, "skolkamrat|NOUN": 1.33, "synfält|NOUN": 1.33, "underlydande|ADJ": 1.33, "frist|NOUN": 1.33, "fyllning|NOUN": 1.32, "förvarna|VERB": 1.32, "stearinljus|NOUN": 1.32, "enhällig|ADJ": 1.31, "insjö|NOUN": 1.31, "ledsaga|VERB": 1.31, "moderskap|NOUN": 1.31, "undantagslöst|ADV": 1.31, "alldaglig|ADJ": 1.29, "avslappning|NOUN": 1.29, "konduktör|NOUN": 1.29, "lågstadium|NOUN": 1.29, "sportig|ADJ": 1.29, "utsändning|NOUN": 1.29, "villighet|NOUN": 1.29, "glans|NOUN": 1.29, "arvinge|NOUN": 1.28, "häfte|NOUN": 1.28, "mejeri|NOUN": 1.28, "chockera|VERB": 1.28, "eskort|NOUN": 1.28, "tabu|NOUN": 1.27, "avdelningschef|NOUN": 1.27, "pilgrimsfärd|NOUN": 1.27, "rättfram|ADJ": 1.27, "slaktare|NOUN": 1.27, "betecknande|ADJ": 1.26, "patologisk|ADJ": 1.26, "multimedia|NOUN": 1.26, "frånskild|ADJ": 1.25, "krämpa|NOUN": 1.25, "långsamhet|NOUN": 1.25, "mätare|NOUN": 1.25, "oljud|NOUN": 1.25, "slitage|NOUN": 1.25, "kommendant|NOUN": 1.25, "hök|NOUN": 1.25, "rugby|NOUN": 1.25, "snöre|NOUN": 1.25, "vidröra|VERB": 1.25, "dån|NOUN": 1.24, "sanitär|ADJ": 1.24, "stekpanna|NOUN": 1.24, "idol|NOUN": 1.23, "luftkonditionering|NOUN": 1.22, "svärson|NOUN": 1.22, "tejp|NOUN": 1.22, "viskning|NOUN": 1.22, "fatal|ADJ": 1.22, "arbetsam|ADJ": 1.21, "korporativ|ADJ": 1.21, "långfristig|ADJ": 1.21, "snarka|VERB": 1.21, "tunna|VERB": 1.21, "ärta|NOUN": 1.21, "kassaskåp|NOUN": 1.2, "fela|VERB": 1.2, "maskulin|ADJ": 1.2, "radie|NOUN": 1.2, "utväxling|NOUN": 1.2, "växellåda|NOUN": 1.2, "ånga|VERB": 1.2, "försyn|NOUN": 1.19, "glidning|NOUN": 1.19, "planlägga|VERB": 1.19, "feminin|ADJ": 1.18, "kodifiera|VERB": 1.18, "poem|NOUN": 1.18, "kompanjon|NOUN": 1.18, "stygg|ADJ": 1.18, "anstöt|NOUN": 1.17, "betyg(s)sätta|VERB": 1.17, "defekt|ADJ": 1.17, "fadd|ADJ": 1.16, "sittning|NOUN": 1.16, "besk|ADJ": 1.15, "rigorös|ADJ": 1.15, "moster|NOUN": 1.15, "gnida|VERB": 1.14, "ordningsföljd|NOUN": 1.14, "ärorik|ADJ": 1.14, "gnistra|VERB": 1.14, "pyjamas|NOUN": 1.14, "bergig|ADJ": 1.13, "fuktighet|NOUN": 1.13, "inkassera|VERB": 1.13, "laglighet|NOUN": 1.13, "statist|NOUN": 1.13, "nobel|ADJ": 1.12, "beväpning|NOUN": 1.12, "gymnasist|NOUN": 1.12, "kolossal|ADJ": 1.12, "stek|NOUN": 1.12, "uppkalla|VERB": 1.12, "försegla|VERB": 1.11, "konsortium|NOUN": 1.11, "acceptans|NOUN": 1.11, "grammatisk|ADJ": 1.11, "strykning|NOUN": 1.11, "kalcium|NOUN": 1.11, "fasta|VERB": 1.1, "tillfälligtvis|ADV": 1.1, "genomgående|ADV": 1.09, "hänförelse|NOUN": 1.09, "spårning|NOUN": 1.09, "systerson|NOUN": 1.09, "gunga|NOUN": 1.08, "ohyra|NOUN": 1.08, "opublicerad|ADJ": 1.08, "idrottsplats|NOUN": 1.08, "elastisk|ADJ": 1.07, "arrest|NOUN": 1.07, "dill|NOUN": 1.07, "vax|NOUN": 1.06, "pose|NOUN": 1.06, "bullrig|ADJ": 1.05, "spröd|ADJ": 1.05, "tidsskrift|NOUN": 1.05, "handfat|NOUN": 1.04, "kork|NOUN": 1.04, "immun|ADJ": 1.04, "inlämna|VERB": 1.04, "projektering|NOUN": 1.03, "regelbundenhet|NOUN": 1.03, "karavan|NOUN": 1.02, "krabba|NOUN": 1.02, "membran|NOUN": 1.02, "antikvitet|NOUN": 1.02, "brant|NOUN": 1.02, "genomträngande|ADJ": 1.02, "kemikalie|NOUN": 1.02, "kultiverad|ADJ": 1.02, "rumslig|ADJ": 1.02, "tråkighet|NOUN": 1.02, "namnteckning|NOUN": 1.01, "personell|ADJ": 1.01, "ungkarl|NOUN": 1.01, "rättfärdigande|NOUN": 1.0, "sammankoppla|VERB": 1.0, "aktivering|NOUN": 0.99, "mellantid|NOUN": 0.99, "motorbåt|NOUN": 0.99, "reglemente|NOUN": 0.99, "decimal|NOUN": 0.99, "mosa|VERB": 0.99, "olivträd|NOUN": 0.98, "anskaffning|NOUN": 0.96, "gradera|VERB": 0.96, "huva|NOUN": 0.96, "lodrät|ADJ": 0.96, "brodera|VERB": 0.95, "socka|NOUN": 0.95, "systerdotter|NOUN": 0.95, "turkos|NOUN": 0.94, "huvudrollsinnehavare|NOUN": 0.94, "kraftlös|ADJ": 0.94, "spann|NOUN": 0.89, "förbittring|NOUN": 0.93, "metallisk|ADJ": 0.93, "repertoar|NOUN": 0.93, "avspänd|ADJ": 0.92, "butiksägare|NOUN": 0.91, "kännare|NOUN": 0.91, "samtalspartner|NOUN": 0.91, "överväldiga|VERB": 0.91, "rea|VERB": 0.91, "böna|VERB": 0.9, "diagnostisk|ADJ": 0.9, "ställ|NOUN": 0.9, "kontingent|NOUN": 0.9, "projektil|NOUN": 0.89, "avtäcka|VERB": 0.89, "iakttagare|NOUN": 0.89, "atmosfärisk|ADJ": 0.88, "borttagning|NOUN": 0.88, "differentiera|VERB": 0.88, "fysiker|NOUN": 0.88, "mygga|NOUN": 0.88, "orange|NOUN": 0.88, "silke|NOUN": 0.88, "troende|NOUN": 0.88, "borste|NOUN": 0.87, "sparv|NOUN": 0.87, "stränghet|NOUN": 0.87, "nittonde|NUM": 0.87, "i övermorgon|ADV": 0.86, "motsägande|ADJ": 0.86, "käring|NOUN": 0.85, "blus|NOUN": 0.84, "kärnpunkt|NOUN": 0.84, "projektera|VERB": 0.84, "utstyrsel|NOUN": 0.84, "laser|NOUN": 0.84, "knippe|NOUN": 0.83, "presidium|NOUN": 0.83, "kvast|NOUN": 0.83, "plommon|NOUN": 0.83, "ägarskap|NOUN": 0.82, "oxe|NOUN": 0.82, "snabbköp|NOUN": 0.82, "tilltugg|NOUN": 0.81, "sned|NOUN": 0.8, "egenartad|ADJ": 0.8, "bulletin|NOUN": 0.79, "högerhand|NOUN": 0.79, "squash|NOUN": 0.79, "stadsbo|NOUN": 0.79, "simmare|NOUN": 0.78, "inkvartering|NOUN": 0.77, "majs|NOUN": 0.77, "visare|NOUN": 0.77, "oupphörlig|ADJ": 0.76, "bönfalla|VERB": 0.75, "dosering|NOUN": 0.75, "studiekamrat|NOUN": 0.75, "tryne|NOUN": 0.75, "ånger|NOUN": 0.75, "kvarlåtenskap|NOUN": 0.75, "körsbär|NOUN": 0.75, "rakning|NOUN": 0.75, "integral|NOUN": 0.74, "klibba|VERB": 0.74, "sparsamhet|NOUN": 0.74, "tunnland|NOUN": 0.74, "formge|VERB": 0.73, "moderlig|ADJ": 0.73, "pina|VERB": 0.73, "undervärdera|VERB": 0.73, "jetplan|NOUN": 0.73, "auktorisera|VERB": 0.72, "korporation|NOUN": 0.72, "saliv|NOUN": 0.72, "strömbrytare|NOUN": 0.72, "kurera|VERB": 0.71, "legering|NOUN": 0.71, "smaklig|ADJ": 0.71, "terroristisk|ADJ": 0.71, "hemgift|NOUN": 0.7, "avvara|VERB": 0.7, "förhandsvisning|NOUN": 0.7, "marmelad|NOUN": 0.7, "trafikpolis|NOUN": 0.7, "kittel|NOUN": 0.69, "bi|ADV": 0.69, "brådska|VERB": 0.69, "reseledare|NOUN": 0.69, "akustik|NOUN": 0.68, "forcerad|ADJ": 0.68, "tidsschema|NOUN": 0.68, "årtusende|NOUN": 0.68, "anträffa|VERB": 0.68, "rutnät|NOUN": 0.68, "försakelse|NOUN": 0.67, "pluton|NOUN": 0.67, "ägarinna|NOUN": 0.67, "överräcka|VERB": 0.67, "jordgubbe|NOUN": 0.66, "sesam|NOUN": 0.66, "artikulera|VERB": 0.66, "aprikos|NOUN": 0.64, "krage|NOUN": 0.64, "reklamera|VERB": 0.64, "tempus|NOUN": 0.64, "upplag|NOUN": 0.64, "tekniker|NOUN": 0.64, "avläsning|NOUN": 0.63, "knall|NOUN": 0.63, "molnig|ADJ": 0.63, "sårande|ADJ": 0.63, "särprägel|NOUN": 0.63, "variabel|ADJ": 0.63, "yrkesman|NOUN": 0.63, "återuppståndelse|NOUN": 0.63, "manöver|NOUN": 0.62, "myr|NOUN": 0.62, "överse|VERB": 0.62, "atletisk|ADJ": 0.61, "skolflicka|NOUN": 0.61, "atlet|NOUN": 0.61, "debitering|NOUN": 0.61, "huslig|ADJ": 0.61, "postlåda|NOUN": 0.61, "millennium|NOUN": 0.61, "valla|NOUN": 0.61, "armbandsur|NOUN": 0.6, "betäckning|NOUN": 0.6, "brorsdotter|NOUN": 0.6, "brutto|ADV": 0.6, "scarf|NOUN": 0.6, "annullering|NOUN": 0.59, "flanera|VERB": 0.59, "läkarvetenskap|NOUN": 0.59, "mittemot (el. mitt emot)|ADV": 0.59, "apparatur|NOUN": 0.58, "fosterbarn|NOUN": 0.58, "förbluffa|VERB": 0.58, "illamående|ADJ": 0.58, "vrist|NOUN": 0.58, "avskedsansökan|NOUN": 0.57, "blyertspenna|NOUN": 0.57, "invändig|ADJ": 0.57, "postulat|NOUN": 0.57, "ytterlig|ADJ": 0.57, "ungdomstid|NOUN": 0.56, "kabin|NOUN": 0.55, "nödhjälp|NOUN": 0.55, "kuriositet|NOUN": 0.54, "pantsätta|VERB": 0.54, "hake|NOUN": 0.54, "renlighet|NOUN": 0.54, "stjälk|NOUN": 0.54, "överlämning|NOUN": 0.53, "olympiad|NOUN": 0.52, "bräde|NOUN": 0.52, "hålighet|NOUN": 0.52, "realisering|NOUN": 0.52, "tariff|NOUN": 0.52, "bindel|NOUN": 0.51, "sockel|NOUN": 0.51, "animering|NOUN": 0.5, "didaktisk|ADJ": 0.5, "doktorsgrad|NOUN": 0.5, "husgeråd|NOUN": 0.5, "klarvaken|ADJ": 0.5, "bullra|VERB": 0.49, "persika|NOUN": 0.49, "svärdotter|NOUN": 0.49, "upprepat|ADV": 0.49, "genomskinlighet|NOUN": 0.48, "sonson|NOUN": 0.48, "stridslysten|ADJ": 0.48, "teatralisk|ADJ": 0.48, "tyngdkraft|NOUN": 0.48, "progression|NOUN": 0.48, "stadgande|NOUN": 0.47, "infarkt|NOUN": 0.47, "upphängning|NOUN": 0.47, "tesked|NOUN": 0.47, "uppdykande|ADJ": 0.47, "måtta|VERB": 0.46, "singularis|NOUN": 0.46, "dotterdotter|NOUN": 0.46, "syskonbarn|NOUN": 0.46, "veterinär|ADJ": 0.46, "baktala|VERB": 0.45, "påskrift|NOUN": 0.45, "slutta|VERB": 0.45, "farmaceutisk|ADJ": 0.44, "innertak|NOUN": 0.44, "knackning|NOUN": 0.44, "koffert|NOUN": 0.44, "monitor|NOUN": 0.44, "simbassäng|NOUN": 0.44, "trettionde|NUM": 0.44, "utvändig|ADJ": 0.44, "brudgum|NOUN": 0.43, "inneslutning|NOUN": 0.43, "genomresa|NOUN": 0.42, "karakteristik|NOUN": 0.42, "mör|ADJ": 0.42, "genomfart|NOUN": 0.41, "kameraman|NOUN": 0.41, "dotterson|NOUN": 0.4, "koefficient|NOUN": 0.4, "vägavgift|NOUN": 0.4, "adjö|NOUN": 0.39, "betjäning|NOUN": 0.39, "periodiskt|ADV": 0.39, "trofé|NOUN": 0.39, "vokal|ADJ": 0.39, "fjäder|NOUN": 0.39, "himmelsblå|ADJ": 0.39, "trådbuss|NOUN": 0.39, "trasa|VERB": 0.38, "födelsemärke|NOUN": 0.37, "hövlighet|NOUN": 0.37, "konvergens|NOUN": 0.37, "sorgsenhet|NOUN": 0.37, "brorson|NOUN": 0.36, "ringklocka|NOUN": 0.36, "vardaglighet|NOUN": 0.36, "berömdhet|NOUN": 0.35, "förutbestämma|VERB": 0.35, "folie|NOUN": 0.34, "kejsardöme|NOUN": 0.34, "käke|NOUN": 0.34, "rymling|NOUN": 0.34, "serum|NOUN": 0.34, "avresa|VERB": 0.33, "elektriker|NOUN": 0.33, "syrsa|NOUN": 0.33, "turkos|ADJ": 0.33, "äggvita|NOUN": 0.33, "hypotekslån|NOUN": 0.32, "invalid|NOUN": 0.32, "månljus|NOUN": 0.32, "transplantera|VERB": 0.32, "tursam|ADJ": 0.32, "kvalificering|NOUN": 0.31, "skolväska|NOUN": 0.31, "utprovning|NOUN": 0.31, "skollov|NOUN": 0.31, "likkista|NOUN": 0.3, "packe|NOUN": 0.3, "svärmor|NOUN": 0.3, "bäcken|NOUN": 0.29, "förbrukare|NOUN": 0.29, "grönska|VERB": 0.29, "modus|NOUN": 0.29, "studenthem|NOUN": 0.29, "mekaniker|NOUN": 0.28, "översida|NOUN": 0.28, "fullbordande|NOUN": 0.27, "undervåning|NOUN": 0.27, "aritmetisk|ADJ": 0.26, "fela|NOUN": 0.26, "frisersalong|NOUN": 0.26, "fönsterbräda|NOUN": 0.26, "cirkelformad|ADJ": 0.25, "kardinal|ADJ": 0.25, "oföränderligt|ADV": 0.25, "regelvidrig|ADJ": 0.25, "skrynkla|VERB": 0.25, "otvivelaktig|ADJ": 0.25, "sondotter|NOUN": 0.25, "ekolog|NOUN": 0.24, "åska|VERB": 0.23, "femtionde|NUM": 0.22, "gravera|VERB": 0.22, "ortopedi|NOUN": 0.22, "tekanna|NOUN": 0.22, "fyrtionde|NUM": 0.22, "konservator|NOUN": 0.22, "hurra|NOUN": 0.06, "inrikes|ADV": 0.21, "maka|VERB": 0.2, "askkopp|NOUN": 0.19, "fästman|NOUN": 0.19, "hyvel|NOUN": 0.19, "straffspark|NOUN": 0.19, "stött|ADJ": 0.19, "subtrahera|VERB": 0.19, "kakelplatta|NOUN": 0.18, "kasus|NOUN": 0.15, "svärfar|NOUN": 0.18, "dossier|NOUN": 0.18, "nolla|VERB": 0.18, "återgälda|VERB": 0.17, "besk|NOUN": 0.17, "bräda|VERB": 0.17, "dyrkan|NOUN": 0.17, "enfamiljshus|NOUN": 0.16, "förkroppsligande|NOUN": 0.16, "violin|NOUN": 0.16, "mottaga|VERB": 0.15, "nittionde|NUM": 0.15, "oregelbundenhet|NOUN": 0.15, "sjukskötare|NOUN": 0.15, "stockning|NOUN": 0.15, "toffel|NOUN": 0.15, "vattenmelon|NOUN": 0.15, "verkställare|NOUN": 0.15, "vårlig|ADJ": 0.15, "metalltråd|NOUN": 0.14, "genetiker|NOUN": 0.13, "sextionde|NUM": 0.13, "timmerstock|NOUN": 0.13, "bjälke|NOUN": 0.12, "excellens|NOUN": 0.12, "läsesal|NOUN": 0.11, "profylax|NOUN": 0.11, "koordinator|NOUN": 0.11, "poängställning|NOUN": 0.11, "docka|VERB": 0.1, "fjärran|NOUN": 0.1, "territorial|ADJ": 0.09, "grafiker|NOUN": 0.08, "undertröja|NOUN": 0.08, "anfallsspelare|NOUN": 0.07, "blotta|NOUN": 0.07, "förfrågan|NOUN": 0.07, "raffinera|VERB": 0.07, "specificitet|NOUN": 0.07, "begeistring|NOUN": 0.06, "bergskam|NOUN": 0.06, "okultiverad|ADJ": 0.06, "skrynkla|NOUN": 0.06, "statistiker|NOUN": 0.06, "syra|VERB": 0.06, "vinäger|NOUN": 0.06, "upphetsa|VERB": 0.05, "författningsenlig|ADJ": 0.04, "kalsong|NOUN": 0.04, "klagan|NOUN": 0.04, "kvitt|NOUN": 0.04, "planta|VERB": 0.04, "toppen|ADJ": 0.04, "tvåsidig|ADJ": 0.04}