Efter
H:K:M:ttz
nådige
resolution
döms
Oluff
till
sin
odels
och
möderne
jord
be:te
8
mälingar
i
Månsgården
.

Allmogen
lovade
sig
vilja
låta
det
till
villig
finnas
efter
sin
förmåga
.

Samtycktes
och
avdömdes
fastebrev
gives
till
Måns
Eriksson
i
Mo
uppå
någon
jord
\
i
Moo
belägen
/
som
han
till
sig
på
sina
stugbarns
vägnar
/
:
och
dem
vid
tiden
till
återlösen
tillbytt
och
köpt
har
.
näml.
Måns
Ersson
bytt
jord
för
jord
(
mz
)
?

Upplästes
den
Kungl.
hovrättens
resolution
daterat
den
4
November
1653
.

Brofogden
Johan
Mickelsson
,
fullmäktige
gjord
å
Moses
Anderssons
vägnar
i
Härnösand
,
kärade
till
Moses
broders
son
Anders
Pehrsson
i
Giäle
,
efter
en
broder
part
i
be:te
Giäle
liggandes
,
den
han
nu
uti
en
lång
tid
brukat
har
,
och
be:te
Moses
varken
för
sin
fäderne
arvsrätt
eller
lott
till
det
ringaste
bekommit
.

Helje
Larsson
i
Åflo
inlade
i
rätten
en
räkning
,
var
med
han
bevisade
sig
ha
efter
wäll:tt
befallningsmans
givna
sedel
utlagt
proviant
till
majorns
wälb:
Petter
Palms
skvadron
för
Hammerdals
tinglag
,
av
åtskilliga
persedlar
,
vilka
är
nu
värderade
till
åtta
och
en
halv
Rd:r
uti
redo
penningar
.

Nils
Olofsson
i
Ås
är
av
Daniel
Mårtensson
på
Åsen
stämd
till
tings
och
sig
då
absenterede
,
sak
fälles
han
till
3
m:r
för
svarlösa
.

Hans
Olufz
gård
i
Ede
,
vilken
här
efter
för
kronogård
om
3
tunnland
utsäde
beräknas
skola
och
Måns
Eriksson
i
Mo
utbetalar
till
arvingar
och
kyrkan
för
1
2
/
3
tl:d
od
18
rd:r
.
30
rd:r
.

Be:te
Jon
bekänner
att
Måns
kom
till
Fyrås
och
krävde
kronans
rest
såsom
ock
stämde
sig
till
tings
.

Till
samma
prov
förordnades
Erik
Nilsson
i
Åsen
,
med
sig
tagandes
fem
andra
tolvmän
,
som
jorden
bese
och
uppmäta
kunna
.

ANNO
1662
den
25
November
hölls
ordinarie
laga
ting
med
allmogen
av
Hammerdals
tinglag
vedervarandes
kronans
befallningsman
ärlig
och
välförståndig
Daniel
Bertilsson
samt
de
tolv
edsvurna
lagrättssmän
.

I
lika
måtto
publicerades
Kungl.
Maij:tz
utgivna
patent
daterat
Stockholm
d
.
28
september
Ao
1661
.

Sakfälls
alltså
förbe:te
Pher
Olufsson
efter
det
3
kap.
köpmål
till
penningar
...
...
12
d:r
för
sitt
förfalskade
gods
,
och
tag
den
åter
värd
som
köpte
,
och
den
flärd
som
sålde
,
som
lag
för
mår
.

Resolverades
denne
sak
således
att
syn
skulle
om
detta
först
rannsaka
,
och
sedan
sin
dom
vinna
.

Dock
där
emot
ha
Ås
byggarna
böxel
brev
utav
fordom
befallningsman
förskaffat
av
Jacob
Chr
.

Blev
slutet
,
Mårthen
Tedt
detta
att
betala
.
3
.

Anno
1664
d
.
26
November
då
laga
ting
hölls
med
allmogen
uti
Hammerdahl
besvärade
sig
Knut
i
Onsala
hur
såsom
Per
Broddesson
i
Öhn
har
sig
sålt
en
oduglig
kvarn
vilken
sedan
såld
är
till
en
man
i
Medelpad
,
den
sig
och
beklagade
över
samma
kvarn
.

Avlade
tolvmännen
sin
ed
,
uti
all
ting
efter
yttersta
förstånd
,
sig
så
handha
,
som
de
för
Gud
och
höga
överheten
kunna
ansvara
;

(
10
)
Framkom
Cisila
Olofsdotter
och
tillkänna
gav
,
huruledes
en
lapp
Skol
Nils
har
berättat
och
i
tal
låtit
komma
,
det
Ingrid
Jonsdotter
i
Gisselås
har
lagt
en
lapp
sig
att
förgöra
,
på
det
att
hon
honom
,
Olof
Olofson
i
Giselås
,
till
man
bekomma
skulle
,
således
avhindra
friemålet
dem
Cisilia
och
Olof
emellan
,
vilket
lappen
Nils
nu
efter
förfrågan
jämte
flera
bevis
sådant
intet
vid
någon
sanning
vara
,
utan
bevittnades
Olof
Olofsson
,
vilken
först
friade
till
Cisilia
och
sedan
till
Ingredh
vara
till
sådant
rop
och
rykte
största
orsaken
.

Dragon
om
sin
målsägar
sak
är
av
rytt
.
förlikat
.

Och
sedan
efter
dessa
penningars
utgörande
,
måste
han
Olof
Thoresson
,
till
överflöd
utstå
och
göra
skjutsfärder
till
Bräcke
.

Vilka
bem:te
4
rd:r
Erich
Staffansson
genast
återgiva
skall
,
alldenstund
han
efter
laga
stämning
till
Lijdt
A:o
1664
ej
komparera
velat
,
och
då
till
dessa
olaga
procedurer
ej
svara
velat
.

(
23
)
Avsades
det
Nils
Andersson
i
Bredgård
skall
betala
Peder
Olofsson
i
Östnår
4½
rd:r
8
sk:r
utan
vidare
uppskov
.

(
28
)
Nils
Andersson
i
Bredgård
pålades
att
svara
Jakob
Jönsson
länsmannen
i
Lit
till
den
1
.
december
nästkommande
vid
tinget
,
om
de
bäverhus
förstörande
han
honom
föreviter
.

(
10
)
Ryttaren
Hans
Johansson
skall
efter
rättens
gottfinnande
flytta
till
hus
hos
sina
andra
bönder
där
så
länge
hos
dem
förbli
,
som
han
hos
Sven
Stensson
i
Ede
,
uti
Andersgården
tillhållit
har
,
vilket
han
genast
efterkomma
skall
.

(
13
)
Per
Stensson
i
Skarpås
uppbjuder
någon
jord
ibid
förste
gång
köpt
av
Olof
Larsson
i
Skottgården
och
Per
Persson
i
Andersgården
för
8
rd:r
1½
ort
.

(
16
)
Lapplandsman
i
Hammerdahls
lappmark
,
Lars
Larsson
tillika
med
Jöns
Andersson
,
Nils
Andersson
,
och
Anders
Clemetsson
som
har
förliden
söndag
fyllt
sig
fulla
med
brännvin
och
Lars
som
har
ropat
och
skrikit
på
kyrkovallen
när
folket
gick
i
kyrkan
;
skall
därför
arbitrateter
straffas
till
40
mk:r
sm:tt
men
de
andra
,
Jönss
,
Nills
och
Anderss
förskonades
med
40
mk:r
sm:tt
till
hopa
,
uppå
Kungl:
May:t
nådiga
behag
dessa
böter
skola
utmätas
och
levereras
till
kyrkan
i
Hammerdahl
och
de
fattiga
.

(
25
)
Måns
Andersson
Spielle
in
för
den
sittande
rätten
skällde
tolvmannen
Anders
Jonsson
i
Ede
för
medhängare
,
hade
fuller
rätten
gått
fog
att
skärpa
,
men
för
hans
fattigdom
förskonades
han
på
Kungl:
May:tz
nådige
behag
med
3
mk:r
sm:tt
efter
43
kap.
tingmåla
b:n
LL
.

(
26
)
Efter
rätten
gottfinnande
avsades
,
att
emedan
som
Jon
Eriksson
i
Fyrås
,
icke
har
något
förord
gjort
när
han
sålde
sitt
hemman
,
att
hans
syster
,
Karin
Eriksdotters
jordepart
för
3
Rd:r
16
sk:r
skulle
ej
inräknas
i
den
40
rd:rs
summa
,
han
för
gården
bekom
,
utan
nu
be:te
3
rd:r
16
s:r
fordrar
av
Anders
Sjulsson
i
Fyrås
;
erkände
rätten
av
intet
värde
,
helst
emedan
Anders
av
Joen
hela
gården
köpte
,
och
detta
klander
då
ej
omtalade
,
för
än
nu
,
utan
Anderz
Siulsson
därför
befrias
.

Hans
Eriksson
i
Grenås
angav
i
rätten
,
ha
förliden
3die
dag
jul
bytt
en
häst
med
Sjul
Persson
i
Hallen
,
uti
goda
mäns
närvaro
,
som
tillika
med
honom
uti
Granåhs
hembjudna
var
,
n:n
Jon
Eriksson
och
Per
Olofsson
i
Görvik
och
Nils
Olofson
i
Gåxsjö
,
vilka
efter
avlagd
ed
,
hand
å
bok
,
betyga
,
att
Siul
uti
deras
närvaro
bytte
med
Hanss
Erichson
häst
,
och
tillbjöd
honom
emellan
3
Rd:r
.

Men
för
Aarååss
ödeböle
gives
av
kyrkoherden
allena
18
öre
s:m:tt
må
det
vid
anfordran
årligen
erläggandes
,
belöper
Summan
av
bägge
ödebölerne
Aaråss
och
Annåhs
1
d:r
12
th:r
sef:r
m:tt
.

Emellertid
utgives
ej
där
på
faste
brev
.

Emedan
som
ej
nekas
,
det
Hemmingh
i
Görvik
har
i
livstiden
lovat
Märit
Stensdotter
äktenskap
,
och
sedermera
uti
sitt
yttersta
testamenterat
henne
tredje
parten
av
lös
örena
som
är
av
hans
avlingegods
;
ty
finner
rätten
det
skäligt
,
att
be:te
testamente
må
ju
hållet
bli
,
därför
må
arvingarna
henne
ovägerligen
tillställa
utan
vidare
besvär
bem:te
tredje
part
av
lösörena
.

När
det
skett
är
,
vill
rätten
lagligen
i
detta
ärendet
sluta
,
om
Oluf
Larsson
har
makt
till
en
oskylld
försälja
gården
före
han
själv
den
lagbjudit
och
fastebrev
där
å
bekommit
har
.

Sockenskrivaren
Olof
Mårtensson
högeligen
sig
besvärade
över
Ströms
tolvmän
,
Anders
Jönsson
i
Strand
,
Per
Broddesson
i
Öhn
,
Olof
Jonsson
i
Tullingsås
och
Per
Danielsson
i
Grelsgård
som
efter
många
påminnelser
icke
har
utfordrat
och
utpantat
1672
års
lagmans
,
häradshövdings
och
tingsgästnings
penningarna
av
råg
finnarna
,
utan
måste
för
dem
utlägga
och
betala
och
intet
assistans
av
dem
njutit
.

Regementskrivaren
Johan
Johansson
sig
besvärade
det
han
efter
H:r
överst
löjtnantens
högvälborne
Lars
Axel
Mörners
order
och
befallning
överskickade
A:o
1671
ifrån
Häggenås
med
Per
Hansson
i
Lorås
sju
Rd:r
i
plåtar
att
igen
lösa
några
dukater
som
stod
i
Looråås
,
hos
Sven
Persson
i
underpant
.

Gör
det
någon
/
och
uppå
föregången
allvarlig
Förmaning
/
sig
icke
rättar
/
vara
/
efter
laga
Rannsakning
och
Dom
/
räknad
för
en
Avfälling
/
miste
sitt
Ämbete
/
och
förvisas
Riket
.

Den
som
och
alldeles
gör
avfall
ifrån
vår
rätta
Religion
,
straffas
lika
så
/
och
njuter
aldrig
något
Arv
/
Rätt
eller
Rättighet
inom
Sveriges
Gränser
.

Ingen
som
av
främmande
Religion
är
/
skall
understå
sig
/
någon
som
bekänner
sig
till
Vår
Lära
/
det
vare
sig
Tjänstefolk
eller
andra
/
att
tubba
/
draga
eller
truga
till
sin
Gudstjänst
;
Utan
tillhålla
sitt
Tjänstefolk
/
som
är
av
Vår
Religion
,
att
flitigt
gå
i
Våra
Kyrkor
.

Åhörarna
skola
och
sin
Gudstjänst
troligen
och
med
Andäktighet
förrätta
/
samt
uti
Böner
/
Lovsånger
/
Guds
Ords
hörande
och
Sakramenternas
bruk
/
visa
ödmjukhet
och
botfärdighet
/
icke
allenast
med
Hjärta
och
Mun
/
utan
och
med
själva
åthävorna
/
till
den
store
Gudens
Tjänst
och
dyrkan
.

Det
som
utur
Kyrkans
Lärare
/
till
Förklaring
andrages
/
bör
ske
med
beskedlighet
och
sparsamhet
/
och
alldeles
komma
överens
med
Guds
Ord
och
den
rätta
Kristliga
läran
.

När
de
röra
några
höga
och
djupsinniga
Lärostycken
/
och
Kätterska
villfarelser
/
måste
sådant
ske
grundligen
och
korteligen
/
med
gott
Förstånd
/
Saktmodighet
och
Försiktighet
;
Och
när
en
eller
annan
Text
ger
dem
anledning
/
till
att
tala
något
om
världsliga
Saker
och
Beställningar
/
så
måste
allt
sådant
ske
med
Beskedlighet
och
Varsamhet
/
utan
Obetänksamhet
och
Förmätenhet
uti
Tal
eller
omdöme
om
de
Saker
/
som
en
del
intet
förstå
/
och
som
LäroÄmbetet
egentligen
intet
angå
;
skolandes
de
som
sig
härutinnan
förgripa
/
och
med
någon
otidighet
och
otjänlighet
på
Predikstolen
framkomma
/
första
gången
med
näpst
och
hårt
Tilltal
anses
/
och
om
de
oftare
där
med
beträdas
/
alldeles
sättas
ifrån
sitt
Ämbete
/
det
de
således
Missbrukat
och
vanvördat
har
.

På
Aposteldagarna
/
hålles
Predikan
i
Stockholm
och
andra
stora
Städer
/
som
här
till
varit
vanligt
;
Men
de
mindre
/
och
på
Landet
/
hålles
allenast
en
Predikan
/
vilken
begynnes
Klockan
Åtta
.

Därefter
sjungs
en
Vers
,
om
den
Helige
Andes
bistånd
;
Och
själva
Predikan
begynnes
med
Morgonbönen
och
Fader
vår
/
utan
något
vidlyftigt
Förtal
.

Uti
Landskyrkorna
/
begynnes
Ottesången
/
om
Jul
Påsk
och
Pingstdagen
/
så
bittida
/
att
den
kan
vara
ändad
vid
pass
Klockan
Åtta
om
Morgonen
/
och
Högpredikan
Middagstiden
.

Om
någon
i
oträngda
mål
och
förfallolös
/
sådant
själv
försummar
/
eller
andra
där
ifrån
hindrar
/
och
icke
med
Kristligt
allvar
/
skyndar
till
detta
förhör
;
Då
skola
Föräldrar
och
Husbönder
/
utgiva
första
gången
vardera
fyra
öre
Silvermynt
för
sig
/
och
för
vart
Barn
och
Legion
två
öre
Silvermynt
/
dem
Sexmännen
/
var
uti
sin
Rote
utfordra
och
till
Kyrkans
behov
upptaga
skola
.

Prästerna
skola
hålla
wissa
längder
på
alla
sina
åhörare
/
Hus
ifrån
Hus
/
Gård
ifrån
Gård
/
och
veta
besked
/
om
deras
framsteg
och
kunskap
uti
deras
Kristendoms
stycken
;
driva
med
flit
där
på
att
Barn
/
Drängar
och
Pijgor
/
lära
läsa
i
Bok
/
och
se
med
egna
ögon
/
vad
Gud
i
sitt
heliga
Ord
bjuder
och
befaller
.

Det
heliga
Dopet
/
skall
alltid
värdeligen
och
Gudeligen
förrättas
i
Kyrkan
/
när
icke
Nödfall
/
eller
andra
skäliga
Orsaker
är
/
som
fordra
att
Barnet
skall
döpas
hemma
:

Döpelsen
måste
och
/
så
vida
möjligt
är
/
ske
på
någon
Söndag
/
Helgdag
eller
Bönestund
/
när
den
Kristliga
Församlingen
är
tillhopa
/
och
kan
samhälleligen
bedja
Gud
för
Barnet
/
och
uppväckas
till
Andakt
och
vördnad
för
detta
Salighets
medlet
.

Döpelsen
skall
med
Guds
Ord
och
rent
obemängt
Vatten
förrättas
/
utav
de
ordinarie
Predikanterna
i
Församlingen
där
Barnen
födda
är
/
helst
av
Kyrkoherden
själv
/
om
han
är
vid
handen
och
oförhindrad
.

Till
Barnmorskor
eller
Jordegummor
/
skola
Gudfruktiga
/
ärliga
/
nyktra
/
och
i
sådana
beställningar
väl
förfarna
Kvinnor
/
antagas
och
förordnas
/
uti
Städerna
av
Magistraten
,
och
på
Landet
av
Kyrkoherden
och
Kyrkans
Föreståndare
och
Sexmän
.

De
Kvinnor
som
har
avlat
Barn
tillhopa
med
sina
Fästmän
/
och
föda
samt
söka
Kyrkogång
/
för
än
vigseln
tillkommer
/
skola
icke
intagas
som
andra
kyska
Barnaföderskor
/
utan
med
ett
särdeles
Bönesätt
/
som
i
Handboken
är
infört
.

Sammaledes
besatta
Människor
/
när
de
det
begära
/
och
igenom
Guds
Nåd
/
är
fria
för
Satans
Anfäktningar
/
bekänna
Jesum
Christum
för
sin
Frälsare
/
och
bedja
Gud
/
om
Syndernas
förlåtelse
/
förstå
deras
Salighets
stycken
/
och
föra
ett
Kristligt
Leverne
;
Men
ingalunda
de
/
som
är
i
sådant
sitt
elände
Ogudaktiga
.

Skulle
han
ändå
icke
vilja
bättra
sig
/
då
ger
Kyrkoherden
/
sin
Biskop
och
Konsistorium
sådant
tillkänna
/
vilka
skola
stämma
Syndaren
in
för
sig
/
och
honom
allvarligen
förmana
/
och
där
han
sig
intet
omvända
vill
/
sätta
honom
/
till
en
bestämd
tid
/
ifrån
den
heliga
Nattvardens
bruk
/
och
andra
Kyrkans
Friheter
/
vilket
kallas
det
mindre
Bann
.

§
.
V
.
Var
den
som
uti
bann
sitter
/
Dödssjuk
/
och
ångrar
sina
Synder
/
begärandes
Herrens
Nattvard
/
så
måste
Själasörjaren
honom
det
icke
förmena
;
Dock
med
förbehåll
/
att
han
skall
stå
uppenbara
Skrift
/
i
fall
han
kommer
till
hälsan
:

Men
dör
den
Bannlyste
i
sin
Obotfärdighet
/
skall
han
icke
av
någon
Präst
/
eller
uti
Kyrkogård
/
begraven
vara
.

Ingen
Präst
skall
/
för
någon
sin
egen
/
eller
sina
Förvanters
och
anhörigas
Sak
skull
/
vad
Namn
den
och
ha
kan
/
avstänga
någon
ifrån
HERRens
Nattvard
:

§
.
I
.
Folket
skall
/
så
väl
uti
Predikningarna
/
som
vid
Barnaläran
/
undervisas
/
om
en
rätt
sannskyldig
Böns
egenskap
/
Kraft
och
nytta
/
samt
förmanas
/
dagligen
att
åkalla
GUd
/
hemma
uti
Husen
/
så
väl
som
Allmänneligen
och
enhälleligen
i
Församlingen
/
att
ha
Böner
/
Förböner
och
Tacksägelse
/
för
alla
Människor
/
Konungar
och
all
Överhet
/
och
bedja
/
om
allt
det
/
som
både
den
timliga
och
eviga
Välfärden
befrämja
/
och
där
emot
/
all
Skada
/
Olycka
och
Bedrövelse
/
avvärja
kan
.

Om
Högtids
och
Helgdagar
.

När
någon
Högtids
Dag
infaller
på
Söndagen
/
avhandlas
alltid
i
Högpredikan
/
Högtidens
Evangelium
,
och
det
som
till
Söndagen
förordnat
är
/
förklaras
i
Aftonsången
/
uti
Städerna
/
och
Fredagen
näst
där
efter
/
på
Landet
:

Men
om
en
Aposteldag
faller
på
Söndagen
/
skall
Söndags
Evangelium
predikas
i
Högpredikan
/
och
Helgdagens
i
Aftonsången
.

Vem
sig
å
Naturens
vägnar
gifta
må
/
eller
intet
.
2
.

Vad
Rättighet
de
Barn
äga
/
till
att
ärva
Fader
/
som
födas
i
fästom
.
7
.

Missbrukar
någon
sitt
Ämbete
/
och
viger
sådana
Personer
tillsammans
/
vilka
icke
lovligt
är
/
att
binda
Äktenskap
/
så
skall
han
/
efter
som
Vårt
/
där
om
utgångna
Plakat
förvår
/
spisas
med
Vatten
och
Bröd
i
Fängelse
/
en
Månad
/
och
sedan
förvisas
Landet
.

Vi
vill
och
/
för
god
Ordning
/
samt
andra
viktiga
skäl
/
Äktenskap
emellan
Syskonbarn
/
så
hädan
efter
/
som
här
till
/
för
Vår
Undersåtar
ha
förbjudit
.

De
som
intet
kunna
råda
sig
/
eller
de
sina
/
skola
i
Tid
/
låta
deras
Själasörjare
förnimma
/
när
de
/
eller
deras
anhöriga
/
vilja
trolovas
/
att
han
må
varna
dem
för
de
hinder
/
som
dem
till
skada
/
av
Skuld
eller
Svågerskap
/
kunna
i
vägen
ligga
;
Och
skall
ingen
trolovas
/
som
icke
kan
Lutheri
Catechismum
,
och
har
begått
HErrens
Nattvard
.

Men
är
Saken
klar
/
och
han
själv
ej
har
något
tvivelsmål
därom
/
då
må
han
utan
förfrågan
/
saklöst
lysa
.

Kvinno
Personer
/
som
låta
lägra
sig
av
deras
Brudgummar
/
förr
BröllopsDagen
/
skall
en
Prästman
/
om
deras
förseende
eljest
är
uppenbart
/
intet
viga
med
annan
Brudeheder
/
än
den
som
Våra
Stadgar
/
eller
vanlig
Plägsed
/
tillåter
.

Sedan
skall
Klaganden
stämma
sin
Vederpart
till
DomKapitlet
,
varest
alla
Äktenskaps
skillnader
ordentligen
bör
ske
.

Vill
den
brottsliga
Parten
/
förfallolös
/
sig
ej
inställa
/
när
han
är
vorden
stämd
/
då
framter
den
Oskyldiga
/
världsliga
Domen
/
var
igenom
den
andra
Sakfälld
är
/
och
då
fortfar
Biskopen
med
skillnaden
/
såsom
uti
en
klar
och
ostridig
Sak
.

Uti
Ältenskapet
tillåts
och
skillnad
/
när
Man
eller
Kvinna
vid
världslig
Rätt
/
så
väl
av
andra
skäl
/
som
egen
bekännelse
/
beprövas
har
/
under
varande
Äktenskap
/
beblandat
sig
med
någon
annan
/
och
Hor
bedrivit
/
och
den
oskyldige
Parten
intet
vill
låta
sig
försona
;
På
vilken
händelse
/
de
av
Biskopen
och
Kapitlet
skola
åtskiljas
/
således
/
att
den
oskyldige
sägs
fri
ifrån
Äktenskaps
Bandet
/
och
får
begiva
sig
i
ett
annat
Giftermål
/
vilket
den
Brottslige
där
emot
skall
förbjudas
/
så
länge
den
Obrottslige
blir
ogift
:

Men
hur
vida
den
samme
sedan
må
gifta
sig
/
eller
ej
/
det
lämnas
till
Konsistoriets
omprövande
.

Utan
att
vi
må
fast
bli
och
vandra
i
det
saliga
Liv
som
Gud
ibland
oss
av
sin
stora
mildhet
upptänt
har
.

Så
är
ock
väl
flera
sådana
nyttiga
stadgar
,
vilka
ock
en
part
för
den
skull
mena
vara
komna
ifrån
Apostlarna
,
såsom
den
,
Att
barn
skola
döpas
,
så
väl
som
gammalt
folk
,
Vilken
Kristlig
Stadga
de
galna
vederdöpare
nu
anfäkta
.

Ty
annat
förstås
icke
med
det
ordet
Besvärja
,
än
bjuda
,
ja
bjuda
med
ett
allvarligt
och
förskräckligt
trug
och
hot
,
vid
Guds
stränga
dom
och
straff
.

Efter
h
.
K
.
M
.
ock
väl
vet
,
huruledes
Kungligt
ämbete
kräver
icke
allenast
det
,
att
h
.
K
.
M
.
skall
ha
vårdnad
och
omsorg
om
världsliga
saker
,
och
sina
undersåtars
timliga
gagn
och
bästa
,
Utan
jämväl
vad
som
hör
till
Gudomlig
ära
,
och
samma
sina
undersåtars
eviga
gagn
och
välfärd
.

Ja
,
där
hon
ordentligt
med
sakerna
vill
gå
till
verket
,
så
måste
hon
visserligen
till
det
allraförsta
söka
Gudomlig
pris
och
ära
,
så
framt
ock
att
det
skall
kunna
något
väl
tillgå
i
det
världsliga
Regementet
.

Den
mig
ärar
,
honom
skall
jag
ära
,
Men
den
mig
föraktar
,
han
skall
komma
på
skam
.
,
För
den
skull
vara
och
de
Konungar
i
Skrifterna
högt
beprisade
som
sig
om
Gudomlig
ära
,
rätta
och
rena
Guds
dyrkan
,
mycket
har
vårda
låtit
,
såsom
Konung
Dauid
,
Ezechias
,
Iosias
,
losaphat
etc.
Men
tvärt
om
,
de
andra
som
den
rätta
och
av
Gud
själv
stictada
Guds
tjänsten
har
nederlagt
,
såsom
Saul
,
eller
ock
de
som
den
samma
rätta
Gudstjänsten
förvandlade
uti
Avguderi
,
såsom
Ierobeam
,
Achab
Älias
,
och
deras
vederlikar
allt
för
många
gjorde
,
de
samma
vara
i
Skrifterna
förfärliga
undsagda
,
såsom
det
sig
och
med
verket
nogsamma
lät
befinna
,
att
de
samt
med
deras
ogudaktiga
undersåtar
hårdeliga
var
straffade
.

Item
,
Allt
det
jag
bjuder
er
skola
ni
hålla
,
Intet
skola
ni
lägga
där
till
,
och
intet
taga
där
ifrån
.

Därför
måste
ock
alla
,
både
de
som
till
Prästämbetet
nu
komna
är
,
och
de
som
där
till
komma
vilja
,
med
allsom
största
flit
överläsa
och
studera
Bibeln
,
att
de
där
utav
må
rättsliga
lära
förstå
grunden
uti
alla
stycken
och
artiklar
,
som
Evangelie
predikan
och
Kristlig
!!
lära
tillhöra
.

Därför
har
ock
vår
Herre
Christus
lärt
,
att
Evangelie
tjänare
skola
både
vara
trogna
och
snälla
,
Trogna
i
det
att
de
rätt
lära
,
och
utan
skrymtan
och
personers
anseende
,
det
som
till
straffandes
är
straffa
.

Där
ock
några
sådana
Legenda
kunde
finnas
,
och
måtte
väl
för
den
skull
av
Predikstolen
föregiven
vara
,
Så
görs
än
då
icke
behov
,
att
hon
alltsammans
förtäljas
,
utan
är
nog
,
att
Predikaren
rör
om
några
stycken
där
uti
,
de
som
är
förnämligast
,
på
det
Lasten
ju
må
behålla
mesta
tiden
i
predikan
.

Men
Episteln
skall
alla
Helgdagar
uti
Städerna
ock
så
predikat
vara
,
Aftonsångs
tid
,
eller
ock
bittida
om
morgonen
,
där
förfall
icke
är
på
färde
,
och
de
är
förhanden
som
det
göra
kunna
.

Vettvillingar
som
buller
göra
,
skola
ock
ledas
ut
.

Och
borde
oss
Kristna
icke
älska
dessa
kyrkohundar
,
både
för
den
skull
,
att
uti
Tiderna
icke
där
igenom
skall
ske
något
hinder
,
såsom
nu
sagt
är
,
så
ock
för
främmande
nationers
förargelse
och
förtal
skull
.

Item
för
den
slemma
art
och
otukt
dem
följer
,
att
de
där
snarast
skämma
och
väta
,
som
bäst
är
tillpyntat
,
både
vid
Altare
och
annorstädes
.

Men
var
ock
förmaningar
icke
hjälpa
vilja
,
så
måste
både
kyrkostraff
och
världsligt
straff
emot
dem
brukat
vara
.

Sammaledes
ock
om
andra
nödtorftiga
stycken
,
om
vilken
tillförne
något
rört
är
.

Och
skall
han
där
om
för
än
han
går
på
Predikstolen
,
av
Klockaren
eller
av
honom
som
slikt
begär
,
skriftligen
eller
muntligen
undervisat
vara
.

Sedan
bedjer
vi
dig
käre
himmelske
Fader
,
för
din
helga
Kristliga
församling
i
hela
världen
,
fria
,
frälsa
och
bevara
henne
för
allt
ont
,
Tag
bort
ifrån
henne
alla
otrogna
Herdar
och
falska
Lärare
,
som
denna
din
klena
Hjord
,
lika
som
glupande
Ulvar
och
rytande
Lejon
jämmerliga
förskingra
och
förhärja
,
utsänd
och
giv
trogna
Herdar
och
rättsinniga
arbetare
i
dina
Säd
.

Därför
vill
vi
nu
det
göra
med
detta
fattiga
barnet
,
som
en
Kristlig
och
broderlig
kärlek
av
oss
kräver
,
nämligen
,
ha
genom
Döpelsen
till
vår
kära
Herre
och
Frälsare
Jesum
Christum
,
bedjandes
av
allt
hjärta
,
att
han
värdigas
det
således
nådeliga
undfå
,
förlåta
ty
alla
synd
och
smittor
,
det
välsigna
,
och
till
tröst
och
styrkelse
med
den
helga
Anda
rikliga
begåva
,
sig
själv
samt
med
Gud
Fader
och
den
helga
Anda
till
pris
,
dessa
fattig
barnen
till
salighet
,
och
sinne
Kristlig
församling
till
hugnad
och
förökelse
,
Amen
.

S
.
Augustini
och
andra
gamla
Lärares
skrivelse
väl
förnimma
kunna
,
dock
så
att
man
här
med
icke
dess
heller
fördömer
de
församlingar
i
främmande
land
,
som
honom
icke
så
bruka
,
och
är
likväl
ens
med
oss
uti
alla
nödtorftiga
och
rätta
trons
artiklar
,
efter
det
är
villkorligt
,
såsom
ock
mycket
annat
(
där
om
tillförne
talat
är
)
vid
Döpelsen
,
varför
vi
honom
i
Nöddop
icke
heller
bruka
eller
bruka
kunna
.

Till
det
tredje
,
att
han
sådant
med
själva
gärningarna
oss
bevisar
,
där
han
så
nådeliga
undfick
denna
barnen
,
tog
dem
upp
i
famnen
,
lade
händerna
på
dem
och
välsignade
dem
.

Om
Syndabot
,
Skriftemål
och
Avlösning
.

Därför
skall
ock
ingen
,
som
har
råkat
åter
falla
i
någon
synd
,
hon
vare
så
stor
som
hon
kan
,
varken
förtvivla
eller
där
uti
bli
,
utan
strax
med
det
allraförsta
omvända
sig
till
Gud
igen
,
med
ett
ångerfullt
hjärta
och
begära
nåd
.
,
Och
skall
man
här
akta
,
att
nu
icke
talas
om
den
bättring
eller
syndabot
som
vi
allesammans
dagligen
för
händer
ha
måste
,
bekännandes
alltid
in
för
Gud
oss
vara
syndare
,
såsom
vi
ock
visserligen
är
,
i
det
vi
icke
så
fullkomliga
håller
hans
helga
bud
som
oss
borde
,
och
måste
för
den
skull
alltid
så
bedja
,
som
vår
käre
HERre
Jesus
Christus
oss
har
lärt
i
Fader
vår
,
nämligen
Förlåt
oss
våra
skulder
etc.
Om
vilket
Profeten
Dauid
i
Psalmen
ock
så
talar
,
där
han
säger
,
Jag
känner
mina
missgärning
,
och
min
synd
är
allstädes
för
mig
.

Item
,
icke
heller
för
än
han
sådana
bedrivna
last
förlovat
och
försvurit
har
.

Och
ändock
det
synes
en
ringa
ting
vara
med
Bann
,
så
har
det
likväl
i
sanningen
mycket
uppå
sig
,
när
där
med
rätt
handlat
var
,
Därför
må
ock
väl
var
och
en
som
i
sanna
sak
är
bannlyst
sig
frukta
,
och
vinnlägga
där
om
,
att
han
utav
sådana
farligt
Bann
må
förlossat
vara
.

Därför
skall
ock
ingen
bannlysas
strax
att
han
har
råkat
falla
i
någon
uppenbara
last
,
utan
man
skall
straffa
honom
såsom
Christus
lär
,
och
försöka
om
han
således
besinnar
sig
,
och
bjuder
bättring
till
.

Detta
är
min
Lekamen
.

Dock
skola
Kyrkoherdarna
ganska
troligen
undervisa
folket
om
dessa
allmänneliga
böner
,
att
de
icke
kunna
vara
fruktsamma
,
eller
förvärva
Gudomlig
hjälp
,
med
mindre
de
ske
av
botfärdiga
människor
,
vilka
deras
synder
känna
,
bekänna
och
överge
,
bättra
deras
leverne
,
och
åkalla
Guds
namn
av
en
rättsinnig
tro
till
Medlaren
Jesum
Christum
,
Så
framt
vi
icke
ville
vänta
de
svaren
av
Gud
,
som
Esaias
om
talar
sägandes
,
Om
ni
än
uträcker
era
händer
,
så
bortgömmer
jag
dock
min
ögon
för
er
,
och
om
ni
än
mycket
bedjer
,
så
hör
jag
er
dock
intet
,
Ty
era
händer
är
fulla
med
blod
etc.
Därför
skall
ock
folket
vara
förmanat
till
bättring
,
och
ju
väl
berättat
i
sakerna
,
att
ingen
kan
vara
en
rätter
bedjare
,
med
mindre
han
först
är
en
god
syndebötare
.

Så
må
ock
än
nu
några
Latinska
sånger
med
ibland
sjungen
vara
,
för
deras
skull
som
det
Latinska
målet
kunna
eller
ock
lära
skola
.
,
Det
skall
icke
heller
någon
bekymra
i
saken
,
att
med
denna
Kyrksång
har
i
förtiden
varit
ett
ganska
stort
missbruk
,
såsom
ock
med
allt
annat
,
Där
man
har
här
av
gjort
,
lika
som
ett
syndoffer
eller
förtjänst
,
till
att
där
igenom
förvärva
nåd
och
syndernas
förlåtelse
,
varför
ock
dessa
tingest
så
är
förökat
,
att
där
med
nu
på
sistone
har
nästan
ingen
måtta
eller
ände
varit
,
Ty
vi
kunna
väl
(
på
Guds
vägnar
)
rätta
sådana
missbruk
genom
ett
Kristligt
förstånd
,
och
sedan
finna
den
måtto
där
med
,
som
efter
vår
och
tidens
lägenhet
kan
vara
bekvämligast
.

Först
skall
man
tillse
,
att
uti
dessa
Tider
ingen
del
sjungen
eller
läst
var
,
den
icke
antingen
är
själva
Skrifternas
uttryckta
ord
,
eller
ock
där
med
så
klarliga
kommer
över
ens
,
att
där
på
kan
ingen
tvivelsmål
vara
,
Med
vilka
man
strax
ogillar
och
förkastar
alla
Homelier
i
Legender
,
Hymner
och
alla
andra
sånger
,
där
något
inmengis
som
sig
med
Skrifterna
icke
fördrar
,
Efter
som
ganska
mycket
sådant
är
för
handen
i
de
gamla
Tideböcker
,
Dock
här
med
icke
förbjudet
det
göra
som
S
.
Paulus
råder
sägandes
,
Prövar
all
ting
,
och
behåller
det
som
gott
är
.

Varför
ock
enär
saken
sig
så
begiva
och
det
kräva
kan
,
må
man
väl
något
avkorta
Psalmer
och
annat
.

Sammaledes
skola
och
Landsprästerna
beflita
sig
där
om
,
att
de
måg
avskaffa
de
okristliga
Minne
,
som
Bönderna
mycket
pläga
bruka
i
deras
gästebod
,
och
komma
dem
till
att
bruka
i
samma
staden
,
några
av
dessa
Svenska
Psalmer
,
Eller
förvandla
samma
Minne
,
så
att
de
draga
över
ens
med
Skrifterna
.

Vad
där
till
hör
,
som
är
täcka
,
böta
och
bygga
,
det
skola
samma
Domkyrkors
Sysslomän
oförsumligen
bestyra
och
uträtta
,
Därför
skall
ock
vara
vid
var
Domkyrka
en
viss
Sysslomansgård
,
uti
vilken
förnämnda
Sysslomän
med
gårdsfolket
må
ha
sin
förvist
.

Item
Heligsmål
,
såsom
seder
är
på
Landsbygderna
.

Så
är
ock
det
Guds
vilja
,
att
de
som
uti
Äktenskapet
stadda
är
,
skola
hålla
sig
troliga
och
renliga
,
så
att
de
icke
förkränkt
med
hordom
och
olovlig
beblandelse
,
Ty
det
är
en
liknelse
och
ett
egentligt
beläte
till
den
kontrakt
och
delaktighet
som
är
emellan
Christum
och
hans
Församling
.

Därför
skall
ock
intet
Äktenskap
bindas
innan
femte
led
,
såsom
seder
har
varit
,
med
mindre
besynnerlig
orsak
kan
vara
på
färde
,
varför
något
må
vara
några
efterlåtit
,
uti
någon
av
de
leder
som
icke
är
förbjudna
uti
den
helga
Skrift
,
och
roten
icke
är
allt
för
när
.

Den
förste
punkt
länder
där
på
Huruledes
Linnert
Jörensson
nu
i
förgångna
höst
1601
Lät
utskriva
till
knektar
de
Rikaste
bönder
,
och
de
fattiga
sattes
för
gårdarna
.

Då
gruvade
sig
var
man
,
sägandes
,
Gud
bättra
oss
då
fattiga
skatte
dragare
,
skulle
vi
således
bli
av
vår
överhet
avvisade
är
befruktandes
att
icke
genom
slikt
blir
Crimen
lesse
Majestatis
etc.
För
vilken
förre
punkts
beskyllning
nämnden
och
menige
häradsmän
med
en
svuren
ed
Linnert
således
ent
skyllade
att
han
varken
var
vållandes
eller
viljandes
,
att
hans
tjänare
detta
skalke
stycke
bevisade
mot
Håckon
Anundssons
son
i
Biedesiö
.

Till
vilken
punkt
nämnden
och
menige
häradsmän
samhälleligen
svarade
,
att
Linnert
Jörensson
ingen
deras
sin
rätt
hade
förkortat
,
och
ingen
fattig
sin
rätt
förvägrat
genom
sin
vederparts
tunga
taske
eller
andra
mutor
.

Vilket
alltså
vara
till
gånget
Suen
klockares
egna
söner
och
deras
farbröder
,
samt
med
nämnden
och
menige
häradsmän
med
en
svuren
ed
bekände
och
vittnade
.

Föregiver
och
Raffuall
i
sina
beskyllningar
om
en
falsk
avkortning
på
98
och
99
års
räkenskap
,
vilken
Linnert
kronan
skulle
ha
för
snillat
.

Genom
vilket
tillfälle
Raffuall
strax
tog
sig
ett
skälms
anslag
före
,
således
,
att
han
drog
ut
samma
natten
och
stämde
till
hopa
vid
pass
14
personer
,
som
skulle
fånga
Linnert
,
och
kom
med
samma
sitt
anhang
tillika
om
morgonen
igen
till
Linnert
,
emedan
han
än
nu
låg
på
sin
säng
,
och
gick
in
till
honom
och
fordrade
honom
upp
till
sig
,
föregivandes
om
några
andra
värv
och
ärenden
han
hade
till
att
tala
och
handla
med
honom
.

Vad
flera
punkter
anlangar
,
som
uti
Raffuals
klago
register
skriftligen
antecknade
är
,
som
röra
dem
själva
och
deras
räkenskap
an
,
det
"
överhemställa
vi
högbetrodde
kammarråd
och
kamrer
till
att
rannsaka
,
efterdet
oss
här
om
ingen
befallning
given
är
och
icke
heller
kunna
,
alldenstund
vi
icke
hade
här
närwarandes
tillstädes
någon
kammar
skrivare
som
deras
räkenskap
kunde
förklara
etc.
Och
efter
det
att
Linnert
Jörensson
uti
all
denne
föreskrivna
Raffuall
Larssons
beskyllningars
punkter
lagligen
har
sig
förklarat
och
för:ne
beskyllningar
med
nämndernas
och
menige
häradsmäns
sannfärdiga
bevis
förlagt
och
således
,
genom
yttersta
rannsaknings
rättmätige
berättning
oss
här
på
tinget
förekom
,
är
befriat
och
skärskottit
bliven
.

Därmed
frågade
han
honom
till
,
var
om
han
sig
så
bekymrade
.

Bonden
svarade
sig
en
underlig
syn
sett
ha
.

Kom
för
rätta
Oluff
i
Hulta
och
klageligen
gav
till
känna
,
att
en
benämnd
Nils
Jonsson
i
Myresboda
i
Nye
Socken
,
inhyses
man
,
hade
stulit
honom
ifrån
i
hans
kvarn
hus
8
skeppor
mjöl
,
med
en
säck
,
men
tjuven
bekänner
,
att
han
tog
en
spann
är
4
skeppor
.

Och
samma
natt
stal
han
från
Birge
i
Hulte
4
skeppor
råg
av
hans
kvarn
hus
,
men
han
bekänner
2
skeppor
råg
.

Och
för
fyra
år
förliden
stal
han
från
Jöns
i
Slätåckra
en
tunna
mjöl
med
säcken
,
det
han
själva
bekänner
.

Kom
för
rätta
Tore
Bengtsson
i
Torgh
i
Huetlanda
socken
och
Brijta
Jonsdåtter
ibidem
,
vilka
samtliga
här
för
rätta
bekänner
,
huruledes
de
var
i
skogen
och
högg
på
ett
träd
som
de
hade
aktat
sig
för
till
krutbrännaren
och
sålt
för
penningar
,
var
och
samma
gången
en
annan
piga
benämnd
Brijta
Mattisedåtter
strax
hos
dem
i
skogen
och
högg
på
ett
annat
träd
,
och
våra
för:116
pigor
broderbarn
,
och
emot
det
träd
ville
falla
som
Tore
Bengtsson
och
Brijta
Jönsedåtter
högg
på
,
varnade
de
Brijta
Mattisedåtter
vidare
,
att
hon
skulle
vakta
sig
,
vilket
hon
icke
gjorde
,
och
där
med
föll
trädet
neder
och
i
hjäl
slog
Brijta
Mattisedåtter
.

Och
efter
denna
föreskrivna
fullmakt
,
som
själva
byttes
brevet
ytterligare
förmäler
,
tingskötte
welb:
Nils
Siöbladh
och
välaktig
Linnert
Jörensson
beskeden
man
Måns
Ståcke
i
Halsnäs
i
Rampnkulla
socken
och
hans
sydskenne
,
nämligen
Oluff
Ståcke
,
hustru
Ingridh
herr
Peders
i
Ååby
och
hustru
Elin
,
Peders
i
Karckningarp
,
för:ne
Lambåsa
på
denne
villkor
och
förord
,
som
föreskrivet
står
.

Ty
avhänder
för:ne
Måns
Stacke
ifrån
sig
sin
broder
och
sina
systrar
samt
deras
arvingar
för:116
deras
rätta
fäders
jord
i
Faderstårp
i
Nye
socken
och
till
ägnar
den
in
under
welb:
Jon
Göstaffsson
,
hans
systrar
,
och
deras
samtliga
efterkommande
arvingar
till
att
nyttja
,
bruka
och
behålla
till
evärdeliga
ägo
etc.
Vilken
Stångfälling
welbe:lte
Linnert
Jörensson
,
på
welbe:lte
välbördig
Jon
Göstaffssons
vägnar
annammade
.

Därför
hemställdes
denna
sak
till
höga
överheten
efter
sitt
nådiga
behag
här
utinnan
göra
och
låta
.

Kom
för
rätta
Eloff
i
Saxhult
och
gav
till
känna
om
en
ko
som
var
för
honom
ihjäl
slagen
,
och
samma
ko
fanns
död
liggandes
inne
på
Ericks
välde
i
Boa
skögle
,
och
därför
hade
Eloff
tvivelsmål
,
att
Erick
skulle
slagit
kon
ihjäl
,
för
vilket
tvivelsmål
för:116
Erick
någon
tid
förliden
utfäste
en
12
månne
ed
.

Kom
för
rätta
en
kvinna
Marriet
Påffualsdater
benämnd
i
Ekelundstårp
i
Huetlanda
socken
,
vilken
bekänner
här
på
häradstinget
att
hon
hade
stulit
ifrån
Per
i
Wglekär
en
stutt
,
vilken
hon
genom
Ingebors
råd
och
tillstyrkan
slaktade
och
förtärade
hemma
till
sitt
,
och
efter
alla
man
här
på
tinget
fällde
bön
för
henne
,
efter
hon
var
en
utfattig
kvinna
,
vart
saken
så
försonat
att
hon
för
samma
stut
skulle
böta
kronan
och
häradshövdingen
en
oxa
.

Men
bonden
undstack
sig
till
skogs
,
så
att
fogden
intet
bekom
hans
tall
.

Vart
och
för:ne
Jon
Skrivare
på
för:ne
sin
systers
vägnar
förenat
och
förlikat
med
S
.
Östens
syster
,
Kirsten
Håkon
Suens
benämnd
,
om
det
arv
för:ne
Kirsten
påtalade
efter
för:ne
sin
S
.
broder
.

Kom
för
rätta
en
gammal
ryttare
Nils
Jonsson
benämnd
i
Brytiarydh
och
Carll
i
Kålleboda
,
vilka
samtliga
hade
var
annan
till
tala
om
ett
vedfä
dem
emellan
någon
tid
för
liden
skett
var
.

Och
han
är
welb:
Hans
Strängs
landbo
.

Till
Träletarp
åldenskog
allena
.

Ty
ett
barn
fanns
uti
Lindåsa
göl
litet
för
midsommar
av
en
dräng
,
benämnd
Anders
Olsson
i
Hulta
,
vilket
var
lagt
i
en
vit
linpåse
och
kastat
i
gölen
,
och
vid
drängen
metade
efter
fisk
,
såg
han
det
vita
på
bottnen
i
gölen
och
rodde
dit
och
drog
upp
påsen
med
en
stång
,
och
när
han
den
upplöste
,
fick
han
se
barnet
och
vart
förskräckt
och
lade
påsen
med
barnet
där
på
marken
och
gick
hem
och
kungjorde
det
sin
fader
,
Oluff
Persson
.

Bekänner
och
uppenbarliga
här
för
rätta
i
nämndens
och
menige
mans
åhöro
,
att
han
utan
all
medgiven
orsak
,
allena
av
ett
argt
och
skälms
uppsåt
,
hade
åstundat
Linnert
Jörenssons
liv
,
är
och
gods
med
dess
yttersta
fördärv
i
grund
att
ombringa
,
som
själva
hans
beskyllningars
punkter
i
bokstaven
ytterligare
utvisa
och
förmäla
,
vilka
alla
sammans
nu
som
tillförne
gick
Rauall
under
ögonen
.

Då
skulle
han
sig
där
om
under
höga
överheten
applicera
.

Kom
för
rätta
en
dräng
Hans
benämnd
i
Skeda
,
som
hade
lägrat
två
pigor
,
Anna
och
Bengta
nämnligen
,
till
vilket
han
icke
nekade
.

Kom
för
rätta
Per
Hemmingsson
i
Erickshister
i
Huetlanda
socken
,
fullmyndig
på
Peer
Olssons
vägnar
i
Biedesiö
i
Myresiö
socken
,
att
tingsköta
Peer
Börjesson
i
Getinge
en
full
fjärding
i
all
den
södra
Biedesiö
gård
för
penningar
50
marker
.

Då
gick
gossen
till
i
förtvivlan
och
tog
ifrån
Carll
i
Höckåsa
ett
par
silver
spännen
om
sex
marker
och
penningar
51
/
2
marker
.

Sammaledes
efter
att
för:ne
Per
Olson
hade
belägrat
för:ne
Kirstin
Månsedoter
emedan
han
var
trolovad
med
Gertrudh
därför
blev
han
fälld
till
penningar
40
mark
.

Här
till
svarade
herr
Karll
,
att
han
intet
vet
utav
de
penningar
,
utan
vad
ägodelar
som
är
efter
lille
Anna
dem
har
han
uppskrivit
,
som
han
vill
hålla
med
sin
svuren
ed
och
med
så
många
män
som
honom
läggs
före
.

Här
på
gavs
sådan
besked
,
att
för:ne
Nils
skall
fly
sin
broder
till
—
städes
till
nästa
ting
om
han
kan
,
var
och
icke
,
skall
då
vidare
här
om
besked
och
ställes
till
kapitlet
,
efter
tvivelsmål
är
,
att
båda
bröderna
har
här
om
lagt
rad
,
på
det
han
skulle
kunna
bli
av
med
henne
.

Där
till
svarar
Karjn
i
Högakull
,
att
för:116
Per
skräddare
var
hennes
mans
målsman
efter
han
var
hans
farbror
,
och
att
Per
Skräddare
skulle
haft
så
mycket
inne
med
sig
,
och
vittnade
Girmundh
i
Knapenöte
,
att
de
talades
vid
där
om
,
dock
visste
han
ingen
viss
besked
om
någon
viss
förlikning
ej
heller
någon
bevis
på
ingen
sida
.

ANNO
1603
Den
8
november
stod
laga
ting
i
Flaga
utav
Steneberga
fjärding
i
kronans
befallningsmans
närvaro
förståndig
Lenart
Jörensons
.
uppbjudningar
.
halva
skatte
gården
i
Slätåker
Brende
Öshult
Embhulte
torp
halva
Kulle
gård
halva
skatte
gården
i
Girmunderydh
Nämnden
Carll
i
Snärle
Jon
Olson
i
Mörisboda
Jon
i
Mörisboda
Sune
i
Solagårdh
Jon
Gunnarson
i
Jdenäs
Lasse
i
Seffseboda
Jon
i
Såndåker
Girmundh
i
Åhnhult
Arffuidh
i
Addaridh
Suen
i
Skurreboda
,
Anundh
i
Skurreboda
,
Oluff
Ståcke
i
Karsnäs
,
Fram
kom
Per
Bengtson
i
Fouglakull
och
lade
ett
tingskötnings
brev
i
rätta
,
som
Lasse
Helgeson
har
utgivit
Anno
97
den
3
december
,
som
lydde
,
att
föreskrivna
Per
och
hans
brorson
Bengt
Jonson
har
bekommit
tingskötning
på
samma
gård
och
givit
släkten
själv
104
lod
,
och
nu
har
Jon
Gunnarson
i
Jdenäs
,
som
är
föreskrivna
Bengt
Jons
barns
morfar
och
målsman
,
sålt
Knut
Biörnson
halva
gården
i
Foglakull
,
som
Bengt
Jonson
har
köpt
och
bekommit
brev
uppå
med
for:ne
fader
broder
.

Dess
för
utan
har
och
för:ne
Per
Bengtson
och
Knut
utgivit
Hemmingh
Kaxa
i
Tånga
och
hans
barn
penningar
24
daler
,
och
uppbjudes
nu
förste
resona
Fram
kom
Girmundh
i
Klacku
och
talade
till
Måns
i
Hester
om
något
barn
arv
,
som
han
hade
inne
med
sig
efter
hans
dotter
barn
.

Item
Jngridh
Östensdoter
och
hennes
son
Måns
Gummeson
talade
till
sin
farbror
Birge
i
Nötebärgh
och
Suen
i
Stocksbärgh
om
den
mansbot
,
som
de
har
uppburit
av
Jon
skräddare
,
för
det
han
slog
hans
fader
ihjäl
.

uppsteg
för
Rätten
Haanss
Larsson
Akademien
utskickade
,
och
accusando
sig
besvärade
över
Olof
i
Myra
Nämndeman
samt
Larss
i
Buddeby
,
vilka
för
några
års
förlopp
hade
synat
några
åker
och
Äng
ifrån
bemälda
Akademien
uti
Storegårdhen
och
lagt
till
ett
Skattehemman
ibidem
där
Anderss
Persson
en
Ryttare
då
åbodde
,
och
nu
hans
hustru
,
efter
bemälda
sin
Mans
Dödliga
för
Riksens
Fiender
,
frånfall
:

Och
efter
Såsom
ingen
då
visste
av
bemälda
½
ortugland
blev
de
av
Nämnden
ändskyllade
och
Haanss
sökte
Lagligen
den
Jorden
brukat
har
,
om
han
gitter
något
där
vinna
,
och
det
efter
föregången
Laglig
stämning
;
eljest
är
Rätten
okunnigt
hur
stort
öretal
är
till
Skattehemmanet
i
bemälda
By
.
7
.

Finns
sedan
något
som
så
illa
medfaret
är
att
han
ingalunda
kan
det
vedertaga
,
så
var
Rätten
förklarandes
sig
på
dem
som
skäligen
bevisas
kunna
höet
genom
försummelse
,
och
vanrykte
och
genom
otidigt
bärgande
fördärvat
ha
,
på
vilka
och
Nämndeman
i
lika
måtto
,
besked
och
underrättelse
veta
skall
;

kom
fram
för
Rätten
Anderss
och
Olof
i
Anderssbo
,
och
kärade
till
Mårthen
i
Stynssbo
,
om
En
ängsmosse
om
16
Sommar
Lass
,
vilken
han
nu
hävdar
,
och
de
genom
Rågång
förmenade
sig
kunna
vinna
till
Anderssbo
.

Och
om
något
över
blir
/
:
ty
bemälda
hustru
och
hennes
man
vore
intet
ringa
Kronan
skyldiga
:
/
skall
hon
sin
Morgongåva
bekomma
.

Vad
hennes
Stugbarn
vid
komma
som
ännu
alla
omyndigha
är
,
vilka
och
bemälda
hemman
Älsarby
,
Såsom
deras
Fädernes
Jord
,
ägande
är
:
vilket
deras
Farbror
Larss
ibidem
som
deras
Målsman
är
till
bruks
/
:
dem
tillhanda
med
tiden
:
/
antagit
har
,
skall
och
sina
brorsbarn
vilka
är
två
bröder
och
tre
Systrar
,
väl
försörja
med
goda
husbönder
;
dem
han
icke
själv
mäktig
är
att
antaga
:
och
de
Jordebrev
som
på
hemmanet
vara
kunna
,
begärde
han
att
uti
Socknens
eller
kyrkans
kista
måtte
inlevereras
,
och
honom
däruppå
bevis
meddelas
.
13
.

kom
för
Rätten
Anderss
Olofzson
i
Wambstadh
och
klagade
till
Mårthen
i
Strömssbo
,
om
21
stång
Järn
som
för
honom
arresterade
är
,
och
Mårthen
har
honom
Järnet
sålt
,
begärandes
därför
att
Mårthen
hans
fångeman
måtte
honom
Järnet
förskaffa
utur
arresten
,
och
han
sedan
utför
saken
med
Arrendatorn
Peter
Roschet
vid
Forssmarck
,
Nu
tillspordes
denne
Mårthen
var
han
Järnet
bekommit
hade
?
han
svarade
sig
det
ha
fått
av
arbets
folket
vid
Österby
,
däremot
uppvisade
bemälde
Peter
Roschet
en
sedel
given
av
Anderss
Erichsson
vid
Österby
,
förmälandes
att
stridige
Järnet
är
intet
Fransos
Järn
som
där
faller
.
/
.
denne
Anders
Erichsson
skall
först
citeras
och
stå
både
Anderss
i
Vambsta
och
Mårthen
i
Strömssbo
till
rätta
,
medan
han
föregivna
Järnet
synat
och
Prövat
har
.
19
.

Då
framsteg
bemälde
Herr
Nillss
,
och
svarade
:
att
enär
bytet
hölls
i
Skärssta
efter
Salig
Erich
Jönsson
,
framkom
bemälde
Mårthen
och
sålde
honom
Oxen
som
Haanss
i
Sund
till
förning
hade
,
där
dock
Herr
Nillss
intet
väl
visste
vilken
oxen
tillhörde
,
och
lovade
honom
4
Tunnor
Råg
som
bemält
är
;
detta
köpet
skedde
uti
Mårthenss
i
Biöringe
Närvaro
,
vilken
vittnade
att
bemälde
Mårthen
bjöd
honom
Oxen
,
för
bemälda
spannmål
,
dagen
därefter
ledde
Mårthen
oxen
i
Präste
gården
,
och
satte
honom
i
Porthelijdrett
,
tillsporde
honom
herr
Nillss
om
bemälda
köp
,
han
svarade
att
köp
bör
gå
fram
,
vilket
skedde
uti
Olofz
i
Stockby
Närvaro
,
vilken
vittnade
så
sant
vara
som
bemält
är
,
att
Mårthen
således
svarade
,
och
att
han
jämte
Mårthen
ledde
oxen
i
Stallet
,
och
tog
sin
kos
Spannmålen
,
flera
vittnen
förmenade
sig
herr
Nillss
kunna
avstad
komma
om
så
behövs
Blev
efter
tidigt
betänkande
avsagt
,
1
att
emedan
herr
Nillss
intet
fulleligen
visste
vilken
Oxen
tillhörde
2
har
han
honom
köpt
med
vinn
och
vittnom
,
varför
skall
köpet
stånda
,
medan
det
Lagligt
är
.

Och
Oloff
Andersson
har
tillstånd
att
söka
sin
broder
Mårthen
,
som
ännu
lever
,
och
utföra
Saken
emot
honom
,
om
han
ohemult
sålt
har
.
22
.

uppsteg
för
Rätten
välbetrodde
Jonas
Bureus
Junior
till
Yla
etc.
påminnandes
Nämnden
om
det
tvistiga
ärendet
som
länge
här
uti
Rätten
hängt
har
,
emellan
hans
Fader
på
den
ena
sidan
,
kärande
,
:
och
Ädel
och
välborne
Jacob
Fårbetz
etc.
på
den
andra
sidan
,
svarande
,
anlangande
två
Sågkvarnar
,
som
bemälde
Fårbetz
har
för
sju
års
tid
sedan
upprätta
låtit
uti
en
Ström
Elgfhorss
benämnd
,
vilken
han
förmenar
med
rätta
lyda
under
Bännebool
;
men
välbetrodde
Bureus
,
samt
Såtterboerne
,
där
han
och
ägande
är
,
har
stadigt
pretenderat
bemälda
Fors
vara
belägen
på
bemälda
Såtterbyess
ägor
,
:

När
Nämnden
när
Synen
hölls
skulle
som
Lag
säger
sig
förklara
,
begärde
Bureus
dilation
för
några
vittnen
skull
som
intet
tillstädes
vore
,
och
om
denna
handel
vetskap
hade
,
det
honom
ej
förvägras
kunde
.

Sedan
har
Thool
Thomasson
uti
Bool
ofta
och
stadigt
vittnat
och
betygat
på
sin
Sotesäng
där
han
ännu
ligger
,
uti
Mårthenss
i
Bloka
,
Anderss
Perssonss
i
Sotter
,
och
Erichz
i
Rekinde
Närvaro
,
sig
på
åtskilliga
tider
ha
hört
,
först
av
sin
Faders
Fader
,
Thool
i
Gärsta
,
Larss
Erichsson
,
och
av
sin
Fader
Thomass
ibidem
att
de
har
sagt
sig
intet
annat
veta
,
än
att
bemälda
Elgfhorss
har
lytt
till
bemälda
Såtter
,
item
har
bemälde
Larss
Erichsson
,
när
om
bemälda
Forss
talat
blev
,
sagt
till
bemälde
Thool
,
om
du
med
tiden
får
höra
att
det
tvistas
om
Strömmen
Elghfårssen
,
så
minns
min
ord
att
han
lyder
till
Såtter
,
på
denne
hans
Edliga
bekännelse
tillbjöd
de
sin
Ed
avlägga
.

kärade
befallningsman
till
Mårthen
Nämndeman
uti
Faringe
Socken
om
fem
tunnor
kyrkotionde
för
året
1634
,
begärandes
veta
vart
de
är
levererade
,
han
svarade
sig
dem
ha
fört
till
Forssmark
den
24
Martij
,
och
befallningsmannen
därpå
kvittensen
levererat
,
han
nekade
där
till
,
ej
heller
hade
Mårthen
därpå
något
vittne
därhos
,
därhos
sade
befallningsman
om
han
bemälda
kvittens
bekommit
hade
är
det
förkommet
.

Dirich
Keijser
appellerade
etc.
dock
ej
å
Lagmans
ting
som
strax
sedan
hölls
,
sitt
vad
fullföljde
.
31
.

Olof
nekade
sig
där
av
veta
,
Per
Jacobsson
svarade
honom
det
måtte
veta
,
medan
hästen
var
så
lång
tid
där
,
att
han
dog
,
där
hos
arbetade
han
på
en
loge
intet
långt
ifrån
huset
där
hästen
var
:

Olof
sköt
skulden
på
en
knekt
som
ute
är
,
vid
namn
Marcus
,
att
han
där
till
orsaken
vara
skall
.

Således
sententierat
och
avdömt
vara
,
så
bekräftas
denna
Dombok
med
härads
Signet
,
till
yttermera
visso
och
bekräftelse
.

Madz
Erichsson
ibidem
om
ett
våg
led
som
Madz
upprätta
borde
vid
sin
kvarn
,
medan
Thomassess
kvarn
måste
ofta
stanna
uti
bakvatten
,
såframt
vågledet
intet
uppsatt
var
:
men
alldenstund
ingendera
Mjölnaren
var
fullmäktig
,
därhos
kunde
för
detta
ej
heller
rätteligen
Prövas
hur
stort
hålldammen
eller
bemälda
vågled
är
angeläget
,
varför
skola
de
bättre
fullmakt
sig
förskaffa
till
lägligare
tid
,
och
då
skall
om
tvistiga
ärendet
Rannsakas
.
39
.

Johan
Nillsson
beropade
sig
på
Peer
Olofzson
i
Haghgåål
som
Skjutet
synat
har
och
huset
:
han
svarade
Erichz
insaga
vara
fåfäng
,
ty
om
icke
hästen
hade
ränt
med
henne
,
hade
hon
intet
trängt
sig
in
uti
ett
sådant
litet
hus
,
vilket
och
Folk
sett
hade
,
eljest
när
Skjutet
sedan
Låg
på
Marken
,
kom
åter
Erichz
häst
och
Bet
det
ändå
illa
:
men
förra
var
Mankan
sönder
bruten
i
dörren
på
huset
,
varav
det
dött
blev
.

Jämväl
har
Larss
Cnutzson
allena
brukat
en
teg
som
genom
Syn
för
elva
år
sedan
vanns
ifrån
Fingarn
och
det
för
bekostnaden
skull
han
på
synen
använde
.
då
blev
och
när
bemälde
under
Lagman
där
var
,
bemälde
Madz
Grijss
halva
Ängs
teg
i
lika
måtto
tilldömt
:
och
vite
satt
,
vilket
föregivs
Larss
Cnutzson
brutit
ha
,
i
det
han
med
våld
allena
tegen
bärgade
.
52
.

Hustru
Charin
svarade
sig
intet
vara
dess
vållande
utan
hennes
häst
som
räddat
blev
och
emot
hennes
vilja
skenade
på
henne
.

Dessa
blev
förlikta
Nämligen
att
bemälda
hustru
Charin
ger
hustru
Elin
10
daler
koppar
mynt
.
54
.

Då
befallde
och
Befallningsmannen
välbetrodde
Class
Classon
alla
grannarna
uti
byn
att
de
broarna
förfärdiga
skola
var
efter
ägo
sina
.

kom
för
Rätten
Olof
Ramunder
,
och
Ratione
officij
anklagade
Bönderna
på
Gränöön
,
som
Ek
huggit
har
till
deras
Båtar
,
och
därför
på
dem
Dom
begärde
:

blev
avsagt
,
att
Peer
i
Gränöö
skall
leverera
hustru
Ingridh
i
Orthale
en
fjärding
Strömming
på
det
köpet
Han
med
hennes
man
gjort
hade
om
en
Sköta
.

kom
för
Rätten
Sigfridh
i
Gåssvijk
,
och
fem
andra
med
honom
uti
Väddeö
Socken
vilkas
sex
Söner
och
Mågar
unga
och
friska
karlar
,
på
Ålands
hav
omkom
,
enär
de
vore
med
Nillss
Mårtensson
Charselio
i
skjutsfärd
åt
Ålandh
.
och
därför
besvärade
de
sig
alla
accusando
utöver
Länssman
Nillss
Erichsson
,
som
honom
utan
Pass
omlagt
har
,
vilket
om
han
hade
Rannsakat
med
flit
,
hade
de
ännu
som
borta
blev
,
varit
vid
livet
,
medan
Charselio
ingen
omläggning
som
de
menade
,
borde
;
Där
till
bemälde
Länsman
svarade
,
att
enär
bemälde
Charselius
anhöll
hos
honom
om
omläggning
har
han
frågat
honom
efter
Passet
,
av
vilket
han
och
en
Kopia
begärde
efter
välborne
Landshövdingens
Befallning
,
Nillss
Mårthensson
svarade
sig
ha
sådant
Pass
som
gäller
till
Land
och
vatten
,
och
sände
honom
en
kopia
ifrån
Gåssvijk
,
och
förra
än
Länsman
fick
den
låta
för
sig
uppläsa
var
han
sin
kos
,
Passet
hade
välborne
Mälchior
von
Falkenbärgh
utgivit
,
vidare
kunde
för
detta
härutinnan
intet
procederas
,
medan
bemälde
Charselius
intet
tillstädes
var
:
utan
allenast
Käranden
häruppå
Bevis
meddelat
till
välborne
Landshövdingens
Resolution
om
bemälda
Pass
.
57
.

kom
för
Rätten
Anderss
Jönsson
i
Biörnhollmen
och
kärade
till
herr
Madz
Johansson
i
Lindrijss
om
tio
daler
silvermynt
,
vilka
han
honom
länt
hade
,
och
begärde
fördenskull
för
detta
sin
betalning
:
gällen
gjordes
för
13
år
sedan
.

Nu
kunde
för
detta
härutinnan
intet
vidare
procederas
,
medan
bemälde
svarande
intet
tillstädes
var
,
Såsom
och
ej
heller
de
vittnen
som
bemälda
hustru
Charin
sig
på
beropade
som
såg
när
Parlamentet
angick
,
här
med
gavs
henne
bevis
där
med
att
söka
Hans
Nåd
Landshövdingen
,
och
anhålla
att
bemälde
Michill
ett
Säkert
Lejde
bekomma
måtte
.
62
.

kom
för
Rätten
Olof
Ramundher
,
och
anklagade
Erich
Erichsson
i
Lindrijss
på
vilkens
ägor
några
Ekar
förbrända
är
uti
ett
Svedje
Land
,
Erich
svarade
hans
Svåger
och
Skytte
under
Skeboo
ha
haft
ett
Svedjeland
,
och
vad
där
skett
var
,
visste
han
intet
,
utan
där
till
må
bemälde
hans
svåger
Jon
i
Sandtorpet
svara
,
han
kunde
intet
Neka
att
några
är
där
emot
hans
vilja
förbrända
,
tre
Ekar
har
Nämnden
funnit
där
alldeles
genom
Svedje
Eld
förbrända
vara
,
därför
Jon
—
40
₥
för
vartdera
böta
skall
,
efter
Riksens
stadgar
,
Oloff
Ramunderss
på
sin
husbondes
vägnar
Ensak
.

Men
om
Ekarna
på
Vredha
och
Yternäss
ägor
skall
vidare
rannsakas
,
och
erfaras
till
vilkens
behov
de
Ekar
huggna
är
,
och
åtskiljas
det
till
Kronans
Behov
hugget
är
,
Sedan
må
Olof
Ramunder
söka
på
andra
orter
och
intet
vidare
så
länge
dröja
i
denna
tigga
Socken
och
med
sina
långsamma
gästningar
fattigha
allmogen
betunga
och
besvära
.
65
.

kom
för
Rätten
hustru
Valborgh
uti
Össby
i
Broo
Socken
och
gav
tillkänna
sig
på
sin
barns
vägnar
,
och
efter
sin
Saligha
Man
Haanss
Hansson
som
för
Riksens
Fiender
bliven
är
,
vara
ägande
till
—
3½
öresland
Jord
uti
bemälda
Össby
,
där
Jönss
Mårthensson
åbor
,
Likväl
tillfogar
bemälde
Jönss
henne
stort
inpass
:
och
därhos
vill
tvinga
henne
ifrån
hemmanet
,
alldeles
:
där
till
Jönss
nekade
;
och
efter
som
han
äger
mera
där
i
gården
som
är
—
5
½
öresland
förmenade
han
sig
genom
lösen
komma
henne
därifrån
,
efter
Såsom
ViceLagmans
Domen
utgiven
av
välborne
Erich
Geeth
utvisar
,
dock
blev
således
för
detta
avskedat
,
att
medan
bemälda
hustru
Valborgz
Man
är
nyligen
som
bemält
är
borta
bliven
,
hennes
barn
omyndigt
,
och
hon
Ensörjande
,
skall
hon
nu
som
tillförende
åtnjuta
,
det
hon
av
hemmanet
innehar
,
till
dess
antingen
hon
bättre
försedd
blir
,
eller
och
barnet
tillväxt
,
dock
Kronans
Rättighet
förbehållen
,
och
vite
till
—
40
₥
sattes
dem
emellan
,
dem
densamma
skall
utan
gensägelse
erlägga
,
som
andra
inpass
tillfogar
,
eller
trätor
förorsakar
:

Vidare
berättade
Nämnden
,
att
den
Domen
bemälde
Lagman
utgivit
hade
skedde
intet
in
Foro
Competenti
,
utan
uti
Väddöö
Socken
,
dit
detta
Häredet
intet
stämt
var
,
mycket
mindre
Nämnden
och
Hustru
Valborgs
Man
som
svaranden
var
och
Saken
angick
.
vilket
blev
annoterat
,
och
henne
efter
hennes
begäran
Bevis
meddelat
.
68
.

blev
vällärde
etc.
Herr
Anderssess
i
Estuna
skrivelse
för
Rätten
uppläst
,
emot
Erich
Jönsson
i
Khubärgha
,
vilken
hade
emot
föregången
Dom
och
eljest
förbud
understått
sig
att
föra
en
bod
ifrån
Qvillunda
hemmanet
det
hans
vyrdighet
äger
:
han
svarade
sig
intet
vara
förbjuden
,
därför
skall
här
om
vidare
rannsakas
,
om
Boden
begärde
han
dilation
,
till
dess
Anderss
i
Håksbodha
,
vilken
hemmanet
förre
åbott
hade
,
kommer
tillstädes
,
med
vilkens
konsens
han
föregiver
sig
Boden
tagit
ha
.
70
.

Sist
vittnade
Anderss
Erichsson
i
Svänsarfva
,
att
han
av
sin
Syster
hustru
Margaretha
i
Skepthamarss
byn
hört
har
,
att
när
Olof
huggen
blev
,
föll
han
vid
öppen
in
till
Hennes
fötter
emot
några
små
Stenar
,
då
kom
en
ung
dräng
och
slog
efter
honom
,
och
råkade
honom
intet
,
men
intet
visste
hon
ehoo
den
var
.

Då
tillspordes
Härads
Nämnd
,
varuppå
de
sig
grundade
,
enär
de
jämte
underlagmannen
dömde
bemälde
Anderss
Nillsson
,
tillika
med
hans
broder
ifrån
livet
,
medan
rannsakat
är
,
att
han
intet
hade
slagit
Olof
Andersson
med
yxhammaren
bak
på
huvudskålen
,
att
hjärnan
skall
och
där
ha
utflutit
,
De
svarade
samtliga
då
sig
uti
hastighet
intet
annat
Pröva
,
eller
142
.
förnimma
kunna
,
än
att
det
slaget
som
Anderss
först
utgav
,
som
han
bekände
drabba
på
Ryggen
,
har
tagit
bak
på
huvudet
som
domen
förmäler
,
och
således
tillika
vara
ett
dödshugg
,
och
det
därför
:
ty
oftabemälde
Nillss
Peersson
begärde
då
in
för
Rätten
,
att
bemälde
båda
hans
Söner
måtte
båda
tillika
svara
till
dråpet
,
vilket
och
Anderss
Nillsson
bejakade
.
för
andras
förbön
skull
som
bjöd
att
han
sin
broder
hjälpa
ville
,
och
alltså
presumerade
de
dem
båda
var
sitt
dödshugg
utgivit
ha
,
:

Då
tillspordes
Nills
Persson
,
varför
han
sådant
gjorde
?
han
svarade
det
ske
av
hans
ringa
förstånd
,
och
enfaldighet
,
menandes
där
med
så
mycket
kunna
uträtta
,
att
bägge
hans
Söner
intet
skola
mista
livet
,
utan
båda
hjälpas
åt
att
böta
,
helst
medan
rätta
målsäganden
har
sin
rätt
på
böter
eftergivit
,
som
domen
utvisar
,
och
alltså
ursäktade
han
både
underlagmannen
och
Nämnden
,
och
bekände
sig
där
till
vara
orsaken
,
honom
till
ingen
ringa
sorg
,
det
han
intet
ihågkom
,
när
han
genom
sin
oförtänkta
begäran
,
sin
Son
uti
stor
vidlyftighet
fört
har
:
vilken
när
han
dömd
blev
gav
sig
strax
på
flykten
,
och
höll
sig
av
vägen
,
till
S
:

M:ttz
nådige
resolution
tillgoda
,
igenlösa
sin
hustrus
rätte
Odel
och
vederlägga
panten
,
Föregiver
att
husen
är
förfallna
och
bortfört
.

Hans
Pehrsson
i
Löffstadh
och
Oluff
Oluffson
i
Ammer
gick
i
löfte
för
Dråparen
.

Sakfälldes
han
för
stämne
till
3
mk:r

Vart
slutit
och
av
Rätten
dömt
,
Efter
det
26
:

Oloff
Oloffson
\
Biutell
/
uppbjuder
halva
…
tunna
Land
\
Seger
Oluffsons
gård
/
uti
Faanbyn
Seger
Oloffson
i
Fanbyn
om
ett
hundrade
tjugo
RD
.
som
de
är
sig
emellan
\
ense
/
om
,
och
blev
så
beslutat
att
Länsman
och
Tolvmän
skulle
rannsaka
hur
många
syster
och
brorparter
där
då
var
uti
Faanbyn
och
om
befinnes
att
Seger
intet
mer
bör
än
sin
brorpart
,
skall
tagas
tillbaka
utav
Seger
\
honom
/
så
mycket
han
övertagit
haf:r
till
dess
riktiga
besked
finns
att
de
andra
hans
bröder
\
och
Syskon
/
äger
med
deras
vilja
och
nöje
utlösa
.

Löp
.
128
mk:r
där
av
tar
Kronan
En
halvpart
löper
64
mk:r
det
övriga
Målsäganden
och
Tobaks
arrendatoren
.

Och
emedan
b:te
Ryttmst
:
den
nedriga
Rätten
ej
Komparera
ville
kunde
Rätten
ingen
dom
i
Saken
falla
\
gångå
/
utan
blev
Remitterat
till
den
Kongl:Håf
Rätten
;
\
Hans
Excell:
Govene:s
ankomst
och
nästkommande
Lands
Ting
.
/
H:r
Befallningsman
tillsporde
om
han
har
låtit
stämma
honom
\
..

Och
har
först
Slagit
Jon
Siulsson
i
Siönäs
med
en
Kniv
i
armen
så
att
han
tolv
veckor
på
säng
ligga
måste
,
den
andra
Olof
Hansson
slagit
i
ryggen
ett
hugg
att
han
och
till
Sängs
legat
har
tre
veckor
.

(
13
.
)
Uppbjuder
förste
gången
Jöns
Joensson
i
Ösiö
Pedher
Jonssonz
anpart
i
Nordhersiö
.

(
5
.
)
Sammaledes
Mattz
Persson
i
Fanbyn
har
olagligen
och
förliden
vinter
städt
en
Piga
Kerstin
från
Hemming
Simonson
,
skall
därför
efter
bem:te
Kap.
plikta
3
mk:r
Även
så
Pehr
Bengtsson
i
Marset
,
har
förliden
Sommar
legat
pigan
Ingebor
Broddesdotter
från
bem:te
Hemming
Simonson
i
Ränswedh
,
Sakfälldes
därför
Per
Bengtsson
efter
för
bem:te
15
Kap.
Bygg:B
.
till
3
mk:r
Sm:tt
Men
Pigorna
Kerstin
Erichsdotter
och
Ingebor
Broddesdotter
,
skola
refundera
och
erlägga
till
Hemming
Simonsson
var
sina
Års
löner
,
som
han
dem
utfäst
har
,
nembl:n
Kerstin
5
ort
och
Ingebohr
6
ort
,
utan
uppskov
,
förmedelst
4
.
punkten
uti
Kungl.
Plakatet
om
legofolks
Stadgande
,
var
med
de
nu
skola
vara
åtskilda

(
34
.
)
Nils
Iffwarsson
uppbjuder
och
,
Faste
Jonssons
i
Rossbohl
Sal
.

(
40
.
)
Olof
Ewertzon
i
Löste
trädde
för
Rätten
,
framvisandes
ett
lagbjudet
och
lagståndet
Köpebrev
,
Daterat
Brattbyn
den
26
Martij
1663
,
med
gode
mäns
underskrift
,
var
med
bevisandes
,
sig
ha
Köpt
av
h
.
Brita
i
Eede
,
och
hennes
Son
Lars
Mårtensson
,
som
barnens
Måhlsman
Hans
Persson
i
Lösta
,
Ett
Tunnland
Jord
i
Eede
,
men
inga
Hus
på
Tomten
för
28
RD:r
samt
alla
dess
tilliggande
lotter
och
lunder
etc.
Så
emedan
ingen
här
på
klandrade
,
ty
utgafs
Faste
brev
.

Fader
,
Nils
Swensson
i
Sidsiöö
har
för
16
år
sedan
,
av
åtskilliga
rätta
Bördemän
köpt
Ett
Tunnland
Jord
,
och
därför
givit
sin
Svägerska
,
h
.
Sigrid
Tohlsdotter
för
hennes
tillfallne
Arvspart
½
tunnland
11
RD:r
och
Olof
Olofsson
i
Stafre
för
1
½
Mäling
givit
6
RD:r
.

Varför
erkände
Rätten
Skäligt
att
Siul
Hermansson
är
berättigat
efter
8
Kap:
Jord
.
b
.

Joen
Person
i
Båsiö
,
uppbjuder
gården
han
åbor
andra
gången
,
sina
Stugbarn
till
återlösen
emot
78
RD:r
.

Swen
Oloffsson
i
Tamnäss
,
Siuhl
i
Miöösiö
,
Oluff
Swänsson
i
Landhsom
Etc
.
uti
Sundziöö
Församling
det
samma
betyga
.
5
.

Ehuru
väl
Trumpetaren
Petter
Olufsson
månde
uppå
Brudflodz
Extra
ordinarie
Ting
d:26
Martij
1670
utlova
,
att
taga
sin
lägerkvinna
Anna
Keelzd:r
till
äkta
,
den
han
haf:r
avlat
barn
med
och
räckte
så
kyrkoherden
H:r
Pehr
Langh
,
som
Rätten
hand
sig
loven
fullborda
;
Men
såsom
Trumpetaren
har
kommit
uti
erfarenhet
att
be:te
Anna
Kelzd:r
\
har
/
beblandat
sig
med
en
annan
Person
,
Näml.
Skräddaren
Hanss
Johansson
på
Frössö
Jemptemarknen
1670
in
Martio
,
några
dagar
för
han
gjorde
handsträckning
med
denna
Anna
Kelzd:r
,
Hanss
Johansson
är
ej
tillstädes
utan
förresten
till
Norige
,
och
Anna
kan
sig
här
från
\
ej
/
unddraga
haft
beblandelse
med
honom
som
hon
sedermera
har
bekänt
för
Trumpetaren
och
nu
detsamma
till
står
,
ty
till
bjöd
sig
Trumpetaren
heller
vilja
utgöra
böterna
för
sig
,
än
taga
Anna
till
äkta
och
sin
äktenskaps
loven
uppsade
,
alldenstund
Anna
ej
bättre
har
sig
ställt
.

H:r
Nilses
Änka
för
3
år
köpt
har
,
och
nu
klandras
av
Rätta
bördeman
,
för
köpet
lagståndet
blev
,
var
över
Resol:des
Att
Anders
Andersson
på
sin
hustrus
wäg:r
är
berättigat
be:te
tunl:d
och
halva
gård
efter
12
.
14
.

Men
H:r
Carl
svarade
,
Kapten
skall
stå
mig
till
Rätt
…
för
Bössan
,
förorsakades
därför
Kapten
stiga
upp
…
gården
efter
bössan
,
och
när
han
dit
upp
kom
,
gick
H:r
Carl
för
åt
i
Stugan
,
och
slog
dörren
igen
,
och
åter
presenterade
sig
i
fönstret
,
fordrandes
honom
att
slåss
m
…
sig
och
hårdragas
,
Svarades
av
Kapten
det
är
icke
Cavalleurs
,
Utan
sådant
tjänar
Skolpojkar
,
har
H:r
Carl
sagt
du
Hundzfott
,
Hundzfott
,
då
H:r
Kapten
har
slagit
H:r
Carl
en
örfil
i
fönstret
,
där
av
H:r
Carl
har
med
de
orden
utbrustit
,
sägandes
,
du
skall
mista
Huvudet
,
du
skall
förvisas
Landet
,
du
skall
böta
till
Kyrkan
,
Hör
du
Hundzfott
,
det
han
intet
längre
kan
tåla
,
utan
H:r
Kapten
begär
H:r
Carl
må
lagligen
plikta
.

Den
30
Januari
1674
Vittnade
efter
avlagd
ed
,
Regement
skrivarens
Johan
Johanssons
dräng
Nils
Olufsson
,
som
förra
Tinget
låg
sjuk
,
Att
han
om
morgonen
stod
på
åkern
och
körde
Trädet
,
har
Pigan
i
gården
gått
efter
honom
och
bett
hemgå
,
vid
det
han
kom
på
gården
,
kom
H:r
CapiteinAnrep
utur
Regement
skrivarens
stuga
och
H:r
Carl
efter
,
H:r
Carl
bad
Kapten
skulle
ingå
och
förlika
sig
med
värden
vilket
han
ej
gjorde
,
Utan
på
gården
slog
Kapten
H:r
Carl
…
slag
med
Spanskrören
,
följdes
så
till
Porten
,
Där
H:r
Carl
åter
…
uti
H:r
Kapten
,
och
ville
ha
honom
tillbaka
,
Men
slets
sig
H:r
Carl
,
När
de
kom
på
åkern
,
fattade
de
varandra
i
håret
,
då
Kapten
ropade
efter
sina
Karlar
att
skilja
åt
,
och
en
av
dem
har
och
tagit
H:r
Carl
i
håret
,
Men
visste
icke
,
vilken
av
dem
var
,
sedan
de
blev
åtskilda
har
H:r
Kapten
slagit
H:r
Carl
med
spansk
rören
3
slag
Ett
över
Kindbenet
,
där
av
han
fick
blånad
,
ett
över
Huvudet
,
och
det
tredje
över
Axeln
,
sedan
har
H:r
upptagit
3
st.
Stenar
och
kastat
efter
,
När
H:r
Kapten
…
i
båten
,
saknade
han
sin
bössa
,
och
gick
därför
själv
femte
tillbaka
upp
i
gården
,
då
H:r
Carl
gick
in
i
stugan
och
Pigan
stängde
dörren
till
,
Men
Nils
var
där
…
Förstugan
,
den
gången
fick
H:r
Kapten
icke
igen
bössan
Därför
sade
Kapten
,
jag
ser
mig
icke
annat
före
än
jag
skall
göra
Hemgång
,
Vilket
Rustmästaren
Swahnbergh
sade
nej
,
det
må
ni
icke
göra
,
har
H:r
Kapten
upplåtit
fönstret
där
H:r
Carl
innan
för
stod
,
och
honom
spottat
i
ansiktet
och
slagit
en
örfil
och
kallat
Hundzfott
,
då
H:r
Carl
svarade
,
du
må
vara
själv
en
Hundzfott
,
där
med
reste
H.r
Kapten
hemåt
.

Pehr
Bengtsson
,
Knut
Keelssons
Svåger
har
observerat
Fatalia
Juris
och
efter
Sveriges
lag
7
Kap:
Jord.b
.

Tolvman
Erich
Önnesson
i
Rind
vittnade
,
att
Kapten
och
Pehr
Andersson
följdes
bägge
till
sig
,
där
Siul
i
Rind
och
var
tillstädes
,
har
Pehr
Andersson
bekänt
för
sig
har
för
sin
nöd
skuld
måste
giva
sig
till
Dragoun
,
där
de
var
andra
handsträckte
.

Manss
broder
,
Keel
Andersson
,
efter
avlagd
ed
refererade
att
han
har
ihjälslagit
ormen
,
vilken
Dragoun
Anders
sedan
har
tagit
på
Lije
Udden
och
lupit
efter
h
.
Märitz
Son
,
då
h
.
Märit
var
vid
pass
ett
St…ke
där
ifrån
,
Alltså
ej
kunde
förstå
,
att
hon
där
av
blev
förskräckt
,
ej
heller
lät
hon
någon
annan
det
förmärka
som
då
tillstädes
var
,
Ej
heller
har
h
.
Märit
för
sig
eller
,
sin
hustru
bekänt
varit
havande
,
som
dock
b
…
tillhopa
uti
en
gård
och
i
nästa
Stuga
,
mycket
mindre
vet
hur
barnet
är
förgånget
,
eller
det
ringaste
haft
någon
Underrättelse
,
Varken
av
henne
själv
eller
någon
annan
.

Länsman
angiver
det
Fänriken
Petter
Wätterströhm
har
andra
gången
belägrat
Konan
Ingebor
Broddesdotter
,
som
är
havande
bliven
Men
ännu
ej
fött
barn
;
Och
emedan
fänriken
är
utkommenderat
bliven
,
ty
uppsköts
till
nästa
laga
Ting
.

Sammaledes
har
då
Sigrid
uppenbarat
sin
Morsyster
,
Elizabet
Larsdotter
i
Äspnäsoch
hans
Stugdotter
Brita
och
alla
ihop
i
Sambsta
…
såväl
fadern
Lars
,
som
Sonen
Lars
Larsson
,
desslikes
Ingebor
i
Hälle
och
Brundfloo
Socken
,
är
Matmoder
i
Blåkulla
och
,
går
där
med
en
Sammets
Rock
;
Sigrid
har
och
,
då
bekänt
för
Pigan
Karin
,
när
hon
bjöd
henne
sin
Ring
,
att
lära
sig
göra
Puken
,
svarat
,
den
är
snart
gjort
,
När
du
klipper
Skägget
och
Sprerlen
av
getterna
och
annat
Raskeri
och
kasta
utom
dörren
,
så
drar
hon
åstad
och
Suger
fä
.
som
H:r
Carls
och
Länsmans
skriftliga
relation
innehåller
.

Tolvman
Herman
Pehrsson
i
Biörnöön
,
Keel
Persson
i
Giällöön
och
Pehr
Andersson
i
Wärwijken
,
som
av
Länsman
Pehr
Andersson
anbefallda
blev
för
2
år
sedan
att
rannsaka
om
den
tjuvnad
Rustmästarens
Pehr
Hemmingssons
hustru
har
bortvisat
,
då
sal
.

Till
detta
kan
Michel
Anderson
ej
undfalla
,
ju
ha
sagt
för
länsman
,
utan
detta
tillstår
,
och
tillbjuder
sig
vilja
bevisa
.

Blev
avskedat
av
Rätten
att
Läns
och
Tolvmän
skola
hålla
en
Sockenstämma
med
första
tillfälle
,
stämmandes
hela
gället
tillsammans
att
hålla
Socken
räkning
om
inbördes
Tunga
och
Skjutsningar
,
på
det
de
en
Jämkning
skulle
sin
emellan
kunna
hålla
och
med
var
annan
likvidera
.

Dato
blev
av
Rätten
avsagt
,
och
slutit
,
det
Kyrkoherden
Ärevyrdig
H:r
Isaac
Alstadius
skall
nyttja
och
bruka
halva
Erich
Önnesons
i
Rindz
Kvarn
till
dess
Pengarna
3
RD:r
blir
Kyrkoherden
restituerade
för
halva
Kvarn
huset
Siuhl
Hermansson
i
Rind
har
sålt
och
Pgr
.
uppburit
.

Pehr
Månssons
hustru
i
Mohlwijken
,
Kerstin
Torkielsdotter
,
som
Anno
1679
den
11
December
förstod
lag
,
sig
själv
tolfte
befria
,
ej
ha
haft
något
olovligen
beställa
med
den
förrymde
Pehr
Swänsson
i
Bräcke
,
som
hon
är
kommen
i
rop
och
rykte
före
,
kunde
nu
inga
Edgärdsmän
framskaffa
,
allenast
sin
egen
man
Pehr
Månsson
begärandes
ytterligare
Dilation
till
nästa
laga
ting
.

B
.
Åtnjuter
halvparten
40
½
RD:r
och
den
andra
halvdelen
bekomma
Systrarna
h
.
Ingiähl
,
Gertrud
och
Sesilla
,
vartdera
13
½
RD:r
bli
40
½
RD:r
.

Den
Kopparkittel
som
1677
års
dom
innehåller
haf:r
Pehr
Andersson
i
Wärwijken
tillika
med
Pehr
Hemmingssons
hustru
h
.
Ingiähl
tagit
i
förlikning
av
sal:
Anders
Hanssons
Änka
,
och
den
samma
fört
till
Swen
Jansson
i
Knytta
för
Penningar
,
den
Pehr
Hemmingson
i
fjol
igenlöste
,
och
till
Änkan
restituerades
.
\
Målsägande
eftergav
sin
Rätt
/
.

Och
bekänner
sig
dels
i
Penningar
och
dels
i
värde
,
fått
,
och
ifrån
sig
levererat
;
Föregivandes
sig
aldrig
å
Pigans
Vägnar
,
varken
något
begärt
eller
Fått
;
Såsom
Peder
Andersson
kan
intet
bevisa
,
Oluf
Penningarna
å
Pigans
Vägnar
av
fordrat
,
varför
kan
Rätten
intet
obligera
Oluf
samma
Penningar
att
Restituera
.

Dock
i
Underdånighet
till
Höglovl.
Kungl.
Hov
Rättens
nådigaste
omdöme
och
Resolution
hemställt
.

Dato
påmindes
om
Kungl:
Maij:ttz
Plakat
och
påbud
och
i
synnerhet
om
Lego
Jons
Stadgan
och
om
de
förrymda
Knektar
och
om
någon
förspörjes
sådant
i
Sinne
ha
och
vilja
fullborda
att
det
må
bli
Vederbörande
kungjort
.

S:r
M:tt
tagit
av
Erich
i
Bohren
,
var
emot
Michell
exciperar
och
berättar
sig
genom
Halfuar
i
Upbyen
dem
avfordra
låtit
och
varken
dem
eller
Saltet
bekommit
och
Halfwar
nu
genom
döden
avgången
är
.

Men
dagen
därefter
förlossade
Gud
henne
igenom
en
stilla
och
salig
död
.

Så
vara
enhälligt
slutet
och
av
gjort
,
intygar
och
attesterar
vi
.

Torparen
Christopher
Olofsson
uti
Älgsiöstufwan
,
gav
ock
tillkänna
,
att
samma
flicka
ifrån
honom
förlidna
Pingstdag
under
Gudstjänsten
bortstulit
1
st.
ost
,
med
några
linnekläder
,
nämligen
1
st.
Servett
,
1
st
Plistinghalsduk
)
1
st
Kammardukshuva
)
och
något
annat
smått
av
mindre
värde
.
§
3
.

Påstående
icke
allenast
,
att
hon
för
detta
,
utan
ock
för
det
hon
sin
tjänst
flera
resor
förlupit
och
strukit
kring
i
socknen
,
måtte
strängeligen
näpst
bli
.
§
7
.

Den
övriga
församlingen
tog
denna
sak
i
Övervägande
,
och
fann
den
vara
av
en
sådan
beskaffenhet
,
att
för
de
många
käromål
,
som
emot
denna
flickan
,
Anna
Jonsdotter
,
blivit
andragna
och
vedergångna
,
målet
borde
vid
laga
Forum
och
till
nästa
höstting
instämmas
;
emedan
slika
och
så
vidlyftiga
mål
,
icke
kunde
komma
under
församlingens
enskilda
avgörande
,
varthän
ock
vederbörande
anvisade
blev
.
§
11
.

A
)
och
till
församlingens
fattiga
1
dr
16
.
/
.
kmt
,
andra
till
varnagel
och
sig
till
förbättring
.

Varpå
modern
,
uti
allas
närvaro
omständligen
frikallade
hustru
Brita
,
och
både
för
Gud
och
människor
vill
draga
skulden
allena
.
§
3
.

Fördenskull
,
och
emedan
Anders
Nilsson
detta
vittnet
på
intet
sätt
jäva
kunde
,
och
i
övrigt
själva
Faktum
vedergånget
och
tillstått
var
,
befanns
han
efter
Högbemälde
Kungl.
Förordningen
de
Anno
1687
har
gjort
sig
brottslig
till
40
dr
smt
böter
,
§
3
.

Så
påtog
sig
Kyrkoherden
,
att
för
Prästgården
allena
4
Bjälkar
framskaffa
.
§
2
.

Församlingen
svarade
:
att
Hemming
aldrig
givit
fattigdel
vore
en
främling
,
samt
orolig
till
sinnes
,
som
med
de
andra
fattiga
icke
särdeles
skulle
förlikas
.

Anders
Swensson
i
Mostorp
,
med
flera
,
begärde
,
att
åldrige
och
avskedade
soldaten
Johan
Påhles
sköterska
,
skulle
för
sitt
omak
,
av
fattigkassan
årligen
njuta
betalning
.

Härjämte
förkunnades
ock
,
att
varest
någon
av
tresko
och
egenvilligt
försummade
slikt
ifrån
sig
i
rättan
tid
framskaffa
,
varigenom
Kyrkoarbetet
,
i
brist
på
spån
,
efter
förslag
och
uträkning
,
kom
att
studsa
skulle
man
vederbörligen
hos
höga
Landshövdinga
Ämbetet
ansökning
göra
om
handräckning
till
arbetets
eftertryckligare
verkställighet
.

Härvid
påmindes
även
församligen
,
att
uti
detta
ärendet
,
endaste
avseendet
borde
vara
,
att
välja
en
sådan
karl
till
klockare
,
som
kunde
informera
de
små
barnen
uti
läsande
vid
kyrkan
,
och
således
även
med
,
om
det
påfordrades
,
undervisa
dem
något
uti
skrivande
.

Som
Lars
Siösten
ifrån
Tyble
anhållit
om
Fattigdels
åtnjutande
,
dock
utan
att
bo
i
Fattighuset
,
ty
äskade
Pastor
Församlingens
utlåtelse
häröver
,
blivandes
honom
hans
åstundan
beviljad
.
§
11
.

Uppräknades
de
resterande
med
Klockpenningarna
,
som
en
del
nu
betalade
,
de
övriga
tillsades
ock
att
inom
14
dagar
betala
i
annan
händelse
tilltar
man
Kronobetjänterna
om
handräckning
.
§
4
.

Stenta
och
Harstorpa
Rotar
köra
fram
gråsten
till
Klockstapeln
och
Kalkugnen
.

Sammansköt
församlingen
,
efter
Hans
Kungl.
Maijtz
nådiga
befallning
,
på
var
Rök
3
.
/
.
kmt
till
Norköpings
Tyska
Kyrka
samt
av
Sätterierna
,
efter
behag
något
mera
,
som
av
Räkningarna
intagas
kan
§
5
.

Församlingen
beklagade
det
att
Vinteråkföret
så
snart
bortgått
,
men
försäkrade
icke
desto
mindre
,
att
både
bjälkar
och
ved
till
rätta
tiden
framskaffa
.
§
5
.

J
.
Dalenius
,
Pastor
)
loci
Carl
Bengtsson
i
Walla
Per
Persson
i
Stenhulta
Kyrkovärdar
.

Frågade
man
församlingens
närvarande
ledamöter
,
vem
de
tyckte
vara
närmast
,
att
bli
antagen
i
fattigstugan
efter
den
avlidna
vansinniga
pigan
Ingrid
?

Även
blev
avslutet
,
att
hustru
Brita
Olofsdotter
i
Nordanås
,
såsom
allmosehjon
utom
fattighuset
skulle
njuta
någon
understöd
.
§
2
.

Nej
så
blev
ock
henne
förövrigt
skriftligt
attest
lämnat
.
§
8
.

Utfäste
sig
ock
församlingens
närvarande
ledamöter
,
att
vilja
låta
hustru
Karin
Larsdotter
i
Wråå
,
uppbära
den
så
kallade
Brudgåvan
uti
norra
Kvarteret
av
Socknen
,
alldenstund
hon
lämnat
till
sin
Svägerska
i
Biörnkällan
,
sin
Rättighet
,
att
uti
Kåhlmårdz
Rootan
i
stället
för
sig
,
brudstad
upphämta
,
som
eljest
hade
ingen
Rätt
sådant
beneficium
njuta
.
§
8
.

Uppsade
sitt
föreståndarskap
för
de
fattiga
Per
Persson
uti
Prästtorp
och
Simon
Larsson
uti
Foglöö
,
och
blev
uti
deras
ställe
antagna
Per
Johansson
i
Stenta
och
Olof
Johansson
i
Tyble
.
§
5
.

Blev
beviljat
,
att
nya
Bänkar
uti
Korgången
,
på
båda
sidor
,
skulle
förfärdigas
,
emedan
Socknen
är
folkrik
,
och
på
Böne
och
Högtidsdagar
,
är
ganska
trångt
om
rum
.
§
10
.

Begärde
Sexmannen
Nils
Hindricsson
i
Dahl
,
så
väl
som
Per
Erichsson
i
Erstorp
dimision
ifrån
SexmansSysslan
,
och
blev
i
deras
ställe
för
Biurstorpa
Roota
,
Anders
Andersson
uti
Trolldahl
och
för
Båltznäsa
Roota
,
Joen
Persson
i
Horssnäs
,
till
Sexmän
förordnade
.

Upplästes
Kladden
på
Kyrkans
inkomst
och
utgift
för
förflutna
året
,
tillika
med
den
avslutade
KyrkoRäkningen
,
med
dess
vederbörliga
verifikationer
,
varemot
ingen
av
Församlingen
hade
att
påminna
.

Saken
blev
,
efter
begäran
,
under
rannsakande
företagen
:
och
sedan
hustru
Maria
offentligen
hade
tillstått
sin
skuld
,
både
beklagandes
sin
stora
dårskap
,
som
ock
begärandes
tillgift
av
församlingen
,
frågade
vad
Satisfaktion
som
Ferengreen
vidare
påstod
?

Sist
av
alltsammans
angav
Pehr
Pehrsson
i
Qwarntorp
,
huruledes
husfolket
hos
Carl
Olofsson
i
Sörgöhlet
,
Olof
Persson
och
dess
hustru
Maria
Jonsdotter
,
i
sitt
äktenskap
ej
kunna
förlikas
,
men
leva
mäkta
illa
i
det
Olof
behåller
och
förvarar
för
sig
det
han
förtjänar
,
utan
att
draga
försorg
för
sin
hustru
och
barn
,
och
hustrun
likaledes
sig
själv
och
barnen
förbehåller
,
det
hon
till
uppehälle
förvärva
kan
,
varav
stor
osämja
,
trätor
,
bitterhet
och
vrede
dem
emellan
uppkommit
.

Pehr
Erichsson
tillstod
,
att
han
varit
vid
Åstufwan
uti
Erich
Christopherssons
frånvaro
,
men
påstod
,
att
Erich
hade
honom
därom
anmodat
,
uti
ett
visst
ärende
:
det
ock
Erich
Christophersson
närvarande
,
besannade
och
bestyrkte
.

Och
som
respektive
domaren
i
orten
låtit
samma
Testamente
,
vilket
i
detta
år
första
resan
nyttjat
fattighuset
uppå
Pastors
begäran
,
enligt
Testamentets
innehåll
,
inflyta
uti
HäradsRätts
Protokollet
,
ty
blev
Extractum
därav
även
uppläst
.
§
4
.

Församlingens
Invånare
påtog
sig
vid
närvarande
sammankomst
,
i
Sommar
att
reparera
ett
stycke
av
Kyrkogårdsringmuren
,
samt
prestera
till
ett
dagsverke
på
matlaget
,
blivande
vid
den
tillförne
antagna
och
gillade
modellen
med
takets
förfärdigande
över
allt
.

Angav
avlidne
och
drunknade
Johan
Christofferssons
änka
,
hustru
Catharina
uti
Mellangärden
Remmeröö
,
hur
hon
befunnit
sig
ha
någorlunda
skäl
att
misstänka
Hustru
Maria
Jonsdtr
uti
Opgården
Sörgölet
,
för
den
säd
,
henne
blivit
av
pörtet
fråntagen
vid
sista
vinterföret
,
och
när
ännu
mannen
stod
på
bår
:
berättandes
,
att
säden
bestått
av
Råg
,
Korn
och
Havre
tillsammans
blandat
till
3
kappar
)
.

Hr
Inspektor
Kralle
påminde
,
att
framlidna
Komminister
Pastor
)
Hr
Jon
Mellins
)
eller
dess
Förfäders
gravsten
på
Kyrkogården
,
skall
vara
något
av
sitt
ställe
skjuten
eller
rubbad
,
vid
det
tillfället
i
sommars
avlidne
Pehr
Olofsson
uti
Skräptorp
blivit
begraven
;
Man
kunde
på
efterfrågan
,
icke
egentligen
få
veta
,
genom
vars
föreställande
sådant
skett
,
men
utlovade
de
närvarande
anhöriga
av
bemälde
Pehr
Olofsson
,
att
med
det
första
sådant
skulle
behörigen
rättat
vara
.
§
19
.

Till
det
sista
sade
Kyrkoherden
;
att
som
han
igenom
Guds
nåd
,
nästan
uti
14
års
tid
,
haft
äran
att
tjäna
uti
Församlingen
och
in
till
denna
stund
på
ingen
Sockenstämma
,
det
ringaste
ord
talat
om
sina
inkomster
och
rättighet
,
varken
större
eller
mindre
,
utan
alltid
dragit
det
kärliga
förtroendet
till
sina
åhörare
,
att
de
självmant
och
rättrådligen
ifrån
sig
måtte
ha
levererat
,
vad
efter
Kungl.
Förordningar
utgå
bör
;
För
vilken
orsak
skuld
ock
aldrig
Sädestionden
på
åkrarna
räknat
blivit
;
Förklarandes
sig
ej
annat
veta
och
vilja
förmoda
,
än
att
alltsammans
rikligt
vore
,
och
därför
även
tackade
Församlingen
behörigen
,
för
den
avlämnade
Tionden
för
innevarande
år
,
allenast
det
påminnandes
,
att
Tionde
av
ärter
,
lin
,
höstråg
etc.
måtte
icke
bli
av
somliga
förglömt
,
som
kan
hända
,
här
till
skett
,
de
rättsinniga
tar
man
undan
;
uppläsandes
till
den
ändan
,
den
1
.
§
av
Kungl.
Förordningen
den
8
Februari
1681
angående
Prästerskapets
uppbörd
av
allmogen
etc.
Församlingen
svarade
;
så
vore
det
aldrig
skett
,
eller
någonsin
därom
talat
.

Så
vara
passerat
,
betyga
av
St.
Malms
Sakristia
1
November
1741
.

Kralle
,
att
Tionde
av
ärter
som
sås
på
trädet
,
ej
kan
betalas
,
som
han
även
förbehöll
sig
,
och
sade
vara
förr
i
Protokollen
influtit
.

Pastor
frågade
ytterligare
,
om
dagsverken
efter
gårdatalet
eller
matlagen
göras
skulle
?

Alldenstund
med
ringningen
efter
Hennes
Kungl.
Maijtt
.
vår
högst
Saliga
)
drottning
kommer
snart
,
efter
Hans
Kungl.
Maijtt
.
nyligen
utkomna
befallning
till
samtliga
Landshövdingarna
,
att
återvändas
alltdärför
blev
fastställt
,
att
med
samma
ringning
ej
skall
,
enär
Påfwelstorpa
Rooten
,
på
vilken
ringningen
nu
står
,
utgången
är
,
uti
en
annan
Roota
begynnas
,
men
kontinueras
uti
samma
Roota
på
innevarande
vecka
,
med
6
Karlar
om
dagen
,
och
det
tills
i
morgon
8
dagar
,
då
med
ringningen
alldeles
slutas
,
enligt
Hans
Kungl.
Maijtt:s
därom
i
dag
å
Predikstolen
publicerade
nådiga
vilja
.
§
8
.

Fann
Församlingen
skäligt
att
bifalla
,
det
Olof
Olofsson
ifrån
Smedstorp
,
hädanefter
såsom
Skräddare
,
jämte
de
andra
,
må
Församlingen
tillhanda
gå
,
till
prov
åtminstone
på
1
år
tills
vidare
,
och
vara
nu
sin
svåger
Olof
Olofsson
i
Karstorp
nu
åter
och
vid
påfordran
,
Socken
Skräddaren
Sven
Svensson
följaktig
;
helst
som
Olof
Olofsson
,
på
tillspörjande
,
tilltrodde
sig
på
gement
vis
samma
syssla
förestå
kunna
.

Som
nu
något
lidit
med
Timringsarbetet
på
Bryggehuset
uti
Prästgården
,
att
nödigt
vara
ville
med
Församlingen
över
)
lägga
,
hur
bekvämligast
detta
arbetet
skulle
innan
instundande
Midsommar
kunna
till
slut
bringas
;
Ty
frågade
man
hur
de
av
Nämndemannen
Nils
Nilsson
projekterade
2
tjog
Nävrar
,
5Va
tolft
Bölning
Bräder
;
samt
800
st.
TakTorv
till
samma
Byggnad
uppå
Församlingen
utdelas
skulle
?

Förkunnandes
Kyrkoherden
,
att
av
Kyrkans
medel
sådant
vara
väl
betalt
,
men
äskade
Församlingens
utlåtande
,
antingen
Kyrkan
skulle
stå
för
sådan
utgift
,
eller
om
Församlingen
ville
honom
slikt
återbetala
?

Men
till
hittelön
av
kyrkans
medel
,
utnämnde
församlingen
åt
murmästaren
Olof
Henningsson
i
Juhlsätter
3
dr
,
samt
åt
Lars
Larsson
uti
St.
Fräntorp
även
3
daler
kmt
.
§
8
.

Föreställandes
därjämte
;
om
icke
församlingen
)
ville
göra
ändring
med
detta
på
sådan
sätt
:
att
den
som
har
barn
att
vistas
hos
;
och
icke
egentligen
)
för
husrum
skuld
,
nödgas
bo
uti
fattigstugan
,
måtte
sig
benöja
med
ett
sådant
underhåll
,
som
gives
till
allmosehjonen
utom
stugan
,
eller
tillhålles
att
flytta
därin
,
om
han
sina
beneficier
behålla
må
?

I
anledning
därav
att
Regements
skrivaren
I
.
Aulin
,
låtit
igenom
Kommissarien
Landeli
,
anmoda
Kyrkoherden
,
att
han
ville
föredraga
Församlingen
bristfälligheten
på
Tjondebode-taket
,
och
att
nödigt
vore
den
samma
måtte
med
det
snaraste
botas
;
blev
ärendet
behörigen
föreställt
.

Uppvisade
Pastor
den
av
Komministern
uti
St.
Jacob
i
Stockholm
,
ärevördige
Herr
Eric
Gerengii
,
i
Koppar
stuckna
Modeller
till
attester
,
som
hädanefter
komma
att
givas
till
dem
,
vilka
flytta
ur
Församlingen
,
enligt
Riksens
Höglovliga
Ständers
Bevillning
på
sista
Riksdag
;
och
emedan
samma
i
koppar
stuckna
Vittnesbörd
,
efter
Plurimum
)
Venerandi
Consistorii
anordning
,
vore
till
96
st
;
redan
på
Prästmötet
i
sistlidne
)
febr
.
månad
,
för
Kyrkans
medel
inlösta
;
Så
beviljades
att
till
Kyrkan
för
vart
Besked
,
hädanefter
erläggas
må
2
å
3
.
/
.
kmt
.
§
8
.

Som
nu
efter
Socken
StugeProtokollets
innehåll
,
pag.
131
.
§
6
det
tillkom
Sandbäcks
Rota
att
votera
på
någon
husfattigs
inskrivande
uti
den
avlidne
åldrige
Smeden
,
Anders
Olofssons
ställe
ifrån
Ändstufwan
;
Så
blev
ock
,
ehuru
både
den
ålderstigne
Eric
Larsson
i
Ändebohl
,
Sven
Larsson
i
Sandwjken
,
Anders
Philipssons
moder
ifrån
)
Hönswjken
,
och
avlidne
Nummer
Soldaten
Kåhrbergs
moder
,
blev
föreslagna
;
den
ålderstigne
änkan
uti
Stetin
enhälleligen
antagen
,
med
det
uttryckliga
förbehåll
,
att
hon
till
fattighuset
inflytta
skulle
.

Uppå
tjänligt
föreställande
,
meddelade
ock
församlingen
av
sina
Fattig
medel
,
3
dr
kmt
till
sjukliga
mönsterskrivaren
Jacob
Lundbom
,
samt
till
den
ålderstigne
Per
Thomasson
ifrån
Hännicketäppan
6
dr
dito
mynt
,
till
någon
understöd
för
sitt
lilla
och
sjukliga
barn
.
§
26
.

Upplästes
Protokollet
som
hållit
vart
på
sistlidne
Valborgsmässosockenstämman
och
blev
vidkänt
.
§
2
.

Berättade
Kyrkoherden
,
att
hur
tid
efter
annan
,
icke
mindre
Församlingen
med
alldeles
nytt
Tak
år
1729
täckte
sina
rum
uti
Prästgårds
större
Byggning
än
hon
samma
år
sina
rum
även
med
nytt
Tak
försett
,
samt
sedermera
både
Församlingens
så
väl
som
sina
eller
Prästgårds
,
reparerat
nu
med
nya
bräder
,
nu
med
Tjärande
,
och
alltsammans
på
egen
bekostnad
till
både
materialer
och
dagsverken
,
det
likväl
bemälda
Tak
är
ändå
nog
otätt
,
och
gör
märklig
skada
,
när
starka
regn
falla
;
Begärandes
att
Församlingen
över
detta
målet
sig
utlåta
behagade
.

Uppvisades
för
Församlingen
den
över
Kyrkomedlen
,
året
om
hållne
Specialen
på
inkomst
och
utgift
,
och
befanns
,
enligt
verifikationerna
vara
till
alla
delar
riktig
,
som
av
KyrkoHuvudRäkningen
närmare
intagas
kan
.
§
8
.

Beslutades
,
att
den
uti
andra
§
omrörda
Summan
för
Prästgårds
byggnad
,
bör
av
Församlingen
inflyta
till
Kyrkan
per
år
,
nämligen
2
daler
i
vita
mynt
av
vart
helt
hemmantal
,
i
4
år
och
vad
som
sedan
brister
,
på
det
femte
året
,
så
att
hela
Summan
på
var
hel
gård
i
5
år
blir
ungefär
9
daler
9
.
/
.
kopparmynt
,
Börandes
första
betalningsterminen
räknas
ifrån
Valborgsmässodag
sistlidne
till
samma
dag
i
tillkommande
år
,
och
så
vidare
samt
att
bemälda
betalning
äntligen
sker
emellan
Jul
och
Matsmässodagen
om
vintertiden
:
emedan
Församlingens
invånare
då
kunna
ha
bästa
tillfället
att
förskaffa
sig
Penningar
.
§
5
.

Men
blev
däröver
denna
resan
ej
något
visst
slut
träffat
.
§
3
.

Upplästes
Specialen
uppå
kyrkans
inkomst
och
utgift
för
sistlidna
år
,
och
befanns
enligt
presenterade
verifikationer
,
alldeles
riktig
vara
.

Sedan
Pastor
nu
som
ofta
tillförne
uti
Församlingens
allmänna
sammankomster
berättat
,
att
längst
för
detta
,
nämligen
redan
uti
avlidne
Salig
)
Herr
Probsten
Espings
tid
höga
landshövdinge-Ämbetet
fastställt
ett
visst
kvantum
uti
mjöl
och
matvaror
i
denna
Församling
att
årligen
utgivas
till
Hospitalet
,
för
vart
helt
hemman
1
lispund
och
5
marker
mjöl
och
5
mkr
kött
,
och
proportionaliter
på
de
mindre
skattlagda
hemmanen
;
beklagade
Kyrkoherden
högeligen
,
att
en
och
annan
av
Församlingens
invånare
är
så
ganska
tröga
med
bemälda
fattigdels
utgivande
,
utnämnde
denna
resan
besynnerligen
Lars
Gustafsson
i
Porten
och
Lars
Persson
uti
Löpsjötorp
,
helst
i
detta
mål
ej
fullgjort
sin
skyldighet
på
två
års
tid
,
ej
heller
framskaffat
någon
ved
till
fattighuset
,
i
mening
att
kunna
med
skäl
denna
innehållna
fattig
delen
förbehålla
sin
gamla
moder
,
som
likväl
är
i
det
stånd
,
att
hon
sig
själv
kan
försörja
,
och
dessutom
vistas
hos
sin
barnlösa
och
någorlunda
sin
utkomst
havande
son
,
bemälde
Lars
Persson
.

Consistorii
cirkulärbrev
det
efter
högvälborne
Herr
Grevens
och
Landshövdingens
gunstige
bifall
ej
några
förordningar
och
Publikationer
skulle
hädanefter
försändas
igenom
Läns
eller
Fjärdingsmannens
anordnande
ifrån
kyrkan
,
där
de
upplästa
är
,
till
en
annan
,
utan
där
förvaras
emedan
slika
Publikationer
och
förordningar
efter
hög
befallning
,
ofta
flera
resor
böra
läsas
.

Pastor
erkände
med
tacksägelse
detta
välborne
Fru
Rosenholms
goda
uppsåt
,
högst
det
Församlingen
till
mycken
nytta
och
prydnad
lända
skulle
då
det
verkställt
blev
.
§
22
.

Presenterades
Förteckningen
,
som
hållen
var
över
de
i
förliden
sommar
,
här
vid
Kyrkan
av
församlingen
gjorda
dagsverken
.
§
4
.

Avslutades
,
att
Johan
Johansson
uti
Stenta
skulle
undfå
av
sina
medintressenter
Sex
daler
kmt
,
för
sin
resa
till
Nykiöping
,
med
en
Supligue
angående
lindrigare
sätt
att
få
(
uttaga
?
)
Kronotionden
av
dem
som
förlidet
år
lidit
missväxt
.
§
8
.

Sporde
Kyrkoherden
Fattighusets
föreståndare
till
om
den
ofärdiga
gubben
Per
Persson
ifrån
Lundsbolstugan
som
på
sista
Valborgsmässo
Sockenstämma
blev
i
fattighuset
intagen
gör
något
buller
i
bland
de
andra
allmosehjonen
.

Löjtnanten
Lidstrand
,
med
allvarsamma
skäl
,
sig
utlät
,
att
det
,
som
i
detta
mål
en
gång
är
avslutat
,
bör
och
skall
stå
fast
,
både
för
skattlagda
och
oskattlagda
emedan
alla
tillkomma
att
vårda
sitt
fattiga
hus
.

Här
på
befordrades
av
Sexmannen
Anders
Simonsson
uti
Nilstorp
;
Skomakaren
ifrån
Simonstorp
församling
Eric
Olofsson
,
som
här
tills
betjänat
Församlingens
invånare
vid
östgöta
gränsen
med
sitt
arbete
,
så
som
på
prov
,
att
nu
vid
Mantalsskrivningen
få
skrivas
för
församlingen
i
bland
de
andra
gärningsmännen
:

Klagades
mycket
över
gamla
Pigan
Brita
ifrån
Koppartorp
för
det
hon
skall
slå
sig
på
lättja
och
ej
vilja
arbeta
hos
dem
som
henne
vid
tillfällen
på
kalla
;
men
därjämte
skall
vara
svår
och
enträgen
med
tiggande
samt
bruka
snatta
;
Brita
framträdde
och
ville
befria
sig
för
denna
beskyllning
;
men
kunde
inte
göra
sig
fri
;
Varför
hon
efter
undfången
varning
,
lovade
ej
mera
i
dessa
mål
vara
någon
besvärlig
,
eller
visa
snålhet
.
§
24
.

Här
på
stannade
församlingen
i
det
slutet
,
att
Kreymans
änka
en
eller
annan
varnings
grad
undergå
skulle
.

Välborna
Herr
Löjtnant
Lidstrand
tillsade
ock
Häradsdomaren
Nils
Nilsson
i
Remna
,
att
han
med
allra
första
måtte
upprätta
Inventarium
,
efter
avlidne
)
Nummer
)
Soldaten
)
Per
Wallman
,
på
det
barnet
,
som
nu
förmedelst
Herr
Löjtnantens
Kristliga
försorg
,
vårdas
hos
Eric
Johansson
i
Qwabben
till
nästa
Michaelij
,
måtte
något
undfå
i
fädernearv
]
,
utav
sin
stugmoder
.
(
§
16
.
)
Behagade
Församlingen
gunstigt
,
på
Kyrkoherdens
föreställande
,
anordna
av
Fattigkassan
,
till
den
eländiga
Munsterskrivaren
Lundbom
,
6
dr
kmt
.
(
§
17
.
)
Erinrade
Herr
Löjtnant
Lidstrand
,
församlingens
invånare
i
gemen
,
att
när
Stamböcker
ankomma
,
som
nu
nyligen
)
skett
för
Hernösands
Kyrka
,
med
var
en
där
till
giva
,
som
behagar
,
samt
så
mycket
han
har
råd
och
ämne
till
.
(
§
18
.
)
Efter
eget
påstående
,
föravskedades
följande
Sexmän
:

Men
som
Per
Nilsson
ej
sedermera
fullbordat
sitt
löfte
,
så
resolverade
Församlingen
att
bemälda
folk
,
med
det
fordeligaste
skola
avlytta
till
en
annan
ort
,
i
avseende
varpå
Sexmannen
i
roten
,
Johan
Johansson
i
Sörgölet
fick
befallning
,
att
å
Församlingens
vägnar
,
sådant
dem
förtyda
.
§
5
.

Alltså
begärde
Pastor
ödmjukt
,
att
Församlingen
nu
täcktes
däröver
sig
utlåta
.

Varest
Erics
Jonsson
ifrån
Båltsnäs
Soldatstuga
,
samt
gamla
Pigan
Anna
Persdotter
ifrån
Qwarnstufwan
,
nu
för
tiden
vistas
!

Angående
den
i
Fattighuset
vistande
flickan
Kierstin
Olofsdotter
,
som
,
oaktat
många
försök
och
prov
,
ännu
icke
kunnat
bli
restituerad
av
sin
sjukdom
,
behagade
Respektive
Herrskapet
på
Erichsberg
,
sig
igenom
Herr
Löjtnant
Lidstrand
gunstigt
förklara
,
att
framledes
vilja
på
några
tjänliga
utvägar
vara
betänkt
,
som
till
bemälda
flickas
hjälp
kunde
sig
lämpa
.
§
8
.

Begärde
Välborne
Herr
Löjtnant
Lidstrand
,
att
komma
i
erfarenhet
,
vilka
vägar
,
utom
den
allmänna
Landsvägen
,
böra
rätteligen
räknas
för
Sockenvägar
?

Så
vara
passerat
,
betyga
på
Församlingens
vägnar
.

J
.
Dalenius
Pär
Pärsson
i
Högen
sexman
.

Kunnande
Eric
Erichson
med
denna
betjäning
,
så
mycket
bättre
komma
ut
,
som
han
redan
fått
hjälp
av
SandwjiksSonen
,
som
för
detta
varit
i
Björckewjk
.
§
6
.

Geringius
till
,
som
årligen
)
är
BrunnsDoktor
vid
Medewi
,
att
denna
fattiga
drängen
,
som
själv
intet
har
något
att
kosta
på
sig
,
kunde
bli
antagen
i
Lasarettet
vid
bemälda
Brun
,
och
där
få
sin
försörjning
.

Högt
ålderstigna
Änkan
,
hustru
Kjerstin
Ersdotter
)
,
som
sitter
i
hus
i
mellangården
)
,
Walla
,
och
har
för
detta
så
länge
hon
förmådde
,
gjort
församlingen
och
dess
Barnaföderskor
mycken
tjänst
,
kommer
att
hädanefter
åtnjuta
samma
förmån
i
Hospitalet
,
som
den
förra
,
dock
begärde
Sexmannen
Lars
Larson
i
St.
Fräntorp
på
hustru
Kjerstins
vägnar
,
att
henne
frihet
lämnas
måtte
,
förbli
i
lilla
stugan
vid
Walla
till
hösten
,
som
henne
icke
kunde
förvägras
,
så
vida
respektive
Herrskapet
på
Ericksberg
sådant
tillåta
vilja
.
§
21
.

Fick
förlov
efter
begäran
,
ifrån
Sexmanssysslan
Olof
Jonson
i
Dahl
,
Lars
Larson
i
Mauritztorp
,
Pehr
Pehrson
i
Erstorp
,
och
Lars
Jonson
i
Ändebohl
;
och
följande
sattes
till
Sexmän
i
deras
ställen
,
nämligen
Jonas
Olson
i
Dahl
för
Bjurstorpa
Rota
,
Nils
Erson
i
Opsala
för
Giersnäsa
Rota
,
Olof
Erson
i
Båldsnäs
för
KjärrBygdaRotan
,
och
Pehr
Arvidson
i
Fäboda
för
Malmsåhs
Rota
.
§
25
.

För
det
andra
frågades
:
om
någon
hade
sig
bekant
att
Mallmberg
,
under
sin
tjänstetid
hos
framlidne
Bryggaren
Hartman
,
har
någon
gång
,
antingen
skrivit
hustrun
till
,
här
i
orten
,
eller
på
annat
sätt
vårdat
hustru
och
barn
?

Det
var
väl
bekant
,
sålänge
Mallmberg
tjänade
för
Kusk
hos
Välborne
Herr
Ryttmästaren
och
Riddaren
David
Hildebrand
,
att
han
henne
då
understödde
understundom
med
litet
underhåll
;
men
det
berättade
flera
:
att
då
de
på
sina
resor
till
Stockholm
,
dels
varit
anmodade
av
hustrun
,
att
fråga
upp
honom
,
dels
såsom
Släktingar
besökt
honom
,
och
föreställt
honom
hur
illa
han
handlade
med
hustru
och
sina
små
barn
;
har
de
alltid
fått
avigt
tal
och
svar
,
jämte
hårda
och
oanständiga
flereslags
utlåtelser
.
§
4
.

Enligt
erhållen
underrättelse
,
skall
nu
ganska
svårt
stå
att
erhållas
Telgsten
ifrån
öland
som
tillförande
varit
projekterat
att
förbättra
Sockenstugegolvet
med
:

NummerSoldaten
Stenbergs
hustru
fick
ock
löfte
på
6
daler
)
kmt
av
fattigkassan
,
för
det
hon
lärt
änkans
i
Västra
Kålberga
Ingrid
Jönsdotter
lilla
dotter
stava
.
§
22
.

Nej
.
4:o
Frågades
om
Barnet
varit
förut
sjukt
?

I
anseende
till
sin
ofärd
ville
väl
Nils
Erson
uti
Opsala
begära
avsked
ifrån
sin
SexmansSyssla
,
som
han
i
2:ne
år
bestridit
hade
;
men
lät
äntligen
övertala
sig
att
vara
Sexman
i
Pålstorpa
Rota
till
hösten
första
gången
.
§
16
.

Sedan
igenom
Respektive
LandshövdingeÄmbetets
remiss
,
under
den
)
11
januari
1757
,
till
överjägmästaren
Winblad
,
Församlingen
erhållit
tillstånd
,
att
,
till
sin
den
tiden
tillärnade
,
nu
fullbordade
,
MagasinsByggnad
,
få
av
Kronans
allmänning
,
Fyrahundra
timmer
,
och
man
åren
tillförne
icke
hunnit
,
att
till
Kyrkan
framskaffa
mera
än
161
.
st.
Stockar
,
så
att
för
Församlingens
räkning
,
ännu
återstå
239
.
dito
,
vilka
på
Kyrkans
bekostnad
,
för
1
år
sedan
,
är
utsynta
och
krönta
,
det
Församlingen
nogsamt
kunnigt
är
;
Fördenskull
och
alldenstund
man
kommit
i
erfarenhet
,
att
en
ny
utsyning
på
Timmer
,
av
krono
allmänningen
skall
snart
ske
,
och
man
således
har
anledning
att
frukta
,
det
Församlingen
torde
komma
att
brista
på
sin
Summa
,
som
vore
en
stor
och
obotlig
skada
,
så
vida
trovärdigt
folk
berätta
,
det
ej
många
parker
på
allmänningen
,
är
med
duglig
skog
försedde
,
så
föreställde
Pastor
,
med
flera
skäl
,
nödvändigheten
,
att
vid
första
vinterföre
,
framskaffa
den
ovannämnda
Summan
.

Gavs
även
tillkänna
,
att
som
Församlingen
på
sista
Mickelsmässo
SockenStämma
,
den
)
16
oktober
sistlidne
,
Se

Begärde
följande
Sexmän
av
sked
;
Nämligen
Sven
Svensson
i
Karstorp
,
som
inemot
20
år
,
haft
denna
Sysslan
:

Och
förordnades
för
Karstorpa
Rota
,
Lars
Olofsson
i
Hällen
,
till
Rotemästare
:

Löjtnant
Anders
Lidstrands
tal
till
Protokollet
uti
SockenStämman
med
Mallms
Socken
,
den
)
1
.

Intet
är
nu
nödigare
att
lappa
,
än
de
revor
som
finnas
på
östra
Gavelns
bägge
hörn
;
vilka
Herr
Ryttmästaren
på
ena
hörnet
nyligen
låtit
emotstödja
;
Men
som
dessa
sprickor
synligen
kommit
av
den
odugliga
grund
,
som
lagd
blivit
till
Kyrkans
skada
,
men
ej
utvidgande
,
och
det
utom
Församlingens
vilja
eller
vetenskap
,
så
påstår
Han
å
Församlingens
vägnar
,
att
den
som
skadan
åstadkommit
,
den
bota
må
,
och
sätta
kyrkan
i
det
stånd
hon
var
,
innan
berörde
odugliga
grund
lagd
blev
.

Ville
Herr
Löjtnanten
gärna
veta
,
om
några
av
de
närvarande
,
kunde
med
säkerhet
säga
:

Men
emedan
ingen
nu
i
hastighet
kunde
härom
tillförlitlig
underrättelse
avgiva
,
blev
målet
till
ett
annat
och
lägligare
tillfälle
uppskjutet
,
då
Herr
Löjtnanten
ville
över
dessa
slags
vägar
Sig
utlåta
.

Utan
skulle
man
endast
söka
till
att
några
andra
små
förbättringar
vid
Kyrkan
göra
,
som
angelägna
vara
kunde
,
såsom
med
Kyrko
och
Torndörrarnas
,
m.m.
stofferande
tillika
med
vad
på
själva
Tornet
kunde
,
till
dess
förvarande
,
nödigt
finnas
.
§
8
.

Upplästes
den
ifrån
Högvördige
Herr
Doktor
och
Biskopen
Jacob
Serenius
till
Kyrkan
ankomne
,
så
kallade
Minneshjälpen
vid
visitationer
,
av
vilken
de
punkter
,
som
kunde
röra
god
ordning
vid
oekonomier
i
Församlingen
)
,
58
)
nu
endast
ventilerades
och
var
följande
,
om
vilka
Församlingen
)
underrättades
.
(
1
)
att
första
Doxologien
näst
efter
Kyrie
läses
ut
helt
och
hållen
,
varest
Kyrie
icke
sjungs
.
(
2
)
Andra
Doxologien
,
näst
för
välsignelsen
,
sker
med
uppstående
av
hela
Församlingen
,
lika
så
för
Trefaldighets
Psalmerna
och
n:o
140
.
(
3
)
Litanian
utelämnas
aldrig
på
Högtids
och
Bönedagar
.
(
4
)
På
SockenStämmorna
uppläses
alltid
3
kap.
Missgärnings
]
balken
)
3
.
4
.
5
.
6
.
7
.
8
.
§§
.
angående
dem
,
som
på
förmaning
sig
icke
bättra
.
(
5
)
Husförhören
skola
börjas
om
hösten
,
sedan
folket
gått
i
tjänsten
.
(
6
)
Vid
årliga
Sockenstämmor
tillsägs
,
att
ingen
som
1
:
a
ggn
vill
träda
i
äktenskap
,
får
vigning
utan
att
kunna
läsa
i
Bok
,
och
Lutheri
Katekes
.
(
7
)
Om
föräldrar
föregå
barnen
med
ond
Exempel
,
sättas
de
ifrån
Herrens
Helige
)
Nattvard
,
och
Tingföras
att
plikta
efter
Missgärnings
)
Balken
)
3
.

Krogar
vid
Kyrkan
upphävas
,
samt
öl
och
brännvins
säljande
vid
gästgiverier
,
för
och
under
Gudstjänsten
,
vid
10
daler
smts
plikt
och
vite
.
(
12
)
Vallgång
av
gossar
förbjuds
,
Se
XI
.

År
1765
den
)
9
Juni
,
kallades
den
närvarande
Församlingen
,
efter
slutad
Gudstjänst
,
in
uti
Sockenstugan
,
då
följande
avhandlades
.
§
1
.

Svarades
enhälligt
nej
.
§
4
.

I
anledning
härav
frågades
:
om
icke
det
vore
billigt
,
att
Kyrkan
för
sina
uti
6
år
utestående
penningar
,
borde
någon
skälig
och
vanlig
Ränta
njuta
?

Jonas
Larsson
uti
Wästergården
,
Remmerö
,
tillika
med
flera
Sockenmän
,
klagade
högeligen
över
den
yppighet
,
som
förövas
av
en
del
unga
drängar
och
gossar
igenom
de
svarta
bandroser
de
tagit
sig
före
att
bruka
uti
halsdukar
med
mera
:
och
kom
Församlingen
enhälligt
överens
,
att
samma
överflöd
och
yppighet
med
det
förra
3
drs
.
vite
,
över
allt
,
för
tjänstedrängar
och
gossar
,
förbjuda
.
§
13
.

Vad
utvägar
borde
vidtagas
,
till
att
ersätta
Fattigkassan
de
utlagde
18
dr
kmt
för
vakthållning
med
mera
,
hos
den
för
detta
sjukliga
Eric
Johansons
hustru
i
Qwabben
,
medan
det
synes
nog
hårt
,
så
vida
mannen
både
bör
och
kunde
sådant
återgälda
,
att
Församlingens
Fattig
Kassa
härmed
må
graveras
?

Vice
Landsmannen
Lars
Samuel
Carell
,
nu
närvarande
,
klagade
högeligen
)
däröver
,
att
Landsvägen
på
Stensjö
backe
,
genom
oaktsamt
sandtagande
i
gropen
,
och
i
kanten
av
vägen
,
blir
alldeles
fördärvad
,
och
är
allaredan
så
mycket
medtagen
,
att
han
snart
stjälper
på
den
ena
sidan
.

Så
tycktes
hans
ord
giva
tillkänna
.

Gud
visste
hur
oskyldig
han
var
,
att
han
var
ohemult
angiven
;
honom
betogs
tillfälle
att
sig
förklara
;
man
ville
honom
nu
fast
oskyldig
,
brottslig
göra
,
med
flera
oanständiga
ord
,
för
vilka
han
behörigen
tilltalades
.
§
5
.

Målet
blev
därför
nu
till
nästa
Söndag
upp
skjutet
för
att
få
de
ovannämnda
vittnen
avhöra
.

Boström
bad
nu
,
i
församlingens
åhöro
,
Jonas
om
tillgift
,
lovade
att
låta
honom
bli
av
sig
oförtalad
,
m.m.
Jonas
eftergav
sin
talan
vidare
,
och
förliktes
med
sin
kontrapart
.

Boströms
Son
Jonas
,
tillstod
icke
allenast
att
han
varit
drucken
,
utan
berättade
även
att
hans
broder
Anders
,
som
tjänar
i
Björkwik
,
hade
givit
honom
brännvin
.

S.D.78
)
uppvisade
bonden
Bengt
Persson
i
Remmerö
och
Soldaten
Nils
Forssberg
,
3
st
nycklar
,
2
av
träd
och
en
gjord
som
en
dyrk
,
dem
Forsberg
tagit
uti
sin
husmans
,
skomakarens
Eric
Perssons
kista
,
under
hans
bortavarande
,
med
utlåtande
,
att
de
hade
skomakaren
misstänkt
för
otrohet
,
så
vida
både
Bengt
och
Forsberg
,
något
saknat
i
sina
hus
,
och
hade
uti
vittnes
övervaro
,
låtit
försöka
besagda
nycklar
,
som
passat
väl
,
den
ena
till
en
Bod
,
den
andra
till
en
loge
i
Remmerö
.
§
2
.

Upplästes
Protokollet
som
hållet
blev
den
17
oktober
sistlidet
år
,
som
till
alla
delar
vidkändes
och
underskrevs
.
§
2
.

Följande
Sexmän
anhöll
om
förlov
:

Februari
innevarande
år
angående
SockenSkolors
inrättande
varöver
Konsistorium
infordrat
Prästerskapets
utlåtande
i
Stiftet
,
m.m.
uti
dess
cirkulär
skrivelse
,
av
den
)
11
.

Församlingens
Ledamöter
fastställde
,
att
alla
de
,
som
låna
penningar
antingen
ur
Kyrkans
eller
de
Fattigas
Kassor
,
böra
hädanefter
erlägga
Intressen
därför
var
gång
MickelmässoSockenstämma
hålls
,
helst
man
trodde
,
att
bättre
tillgång
kan
givas
på
penningar
om
hösten
,
än
om
vårtiden
.
§
6
.

Men
som
pantsilvret
bestående
av
3:ne
silverkoppar
,
1783
uti
augusti
månad
blivit
bortstulna
,
så
frågade
Pastor
församl
:
n
vad
utvägar
skulle
tagas
,
för
att
hålla
både
Kassan
och
låntagare
skadelösa
?

Pastor
lät
församl
:
n
veta
,
att
han
,
i
kyrkovärdarnas
och
fattigföreståndares
närvaro
,
räknat
de
kontanta
penningar
i
Kassorna
och
funnit
dem
vara
alldeles
efter
de
nu
upplästa
räkningarna
,
så
att
Nådårs
Predikanten
)
Mag:r
Herr
redric
Tiselius
redeligen
förvaltat
och
från
sig
lämnat
Kassorna
,
varför
Pastor
å
församlingens
vägnar
honom
betackade
.
§
10
.

Det
berättas
,
att
Orgelverket
,
efter
dess
uppsättande
,
aldrig
blivit
rengjort
,
och
därför
frågade
Pastor
,
om
icke
församl
:
n
ville
anmoda
Herr
OrgelByggaren
,
som
kommer
till
Västra
Vingåker
i
sommar
,
att
rengöra
detsamma
,
samt
,
om
sig
göra
låter
,
att
även
göra
de
stämmor
lindrigare
,
som
nu
tyckas
vara
för
stränga
och
starka
,
i
anseende
till
kyrkan
?
vilket
blev
lovat
.
§
16
.

Pastor
anmälde
,
att
i
anseende
till
den
stora
bristen
på
brödfödan
för
den
arbetande
menigheten
i
Socknen
,
har
församlingens
Patron
Välborne
Herr
Ryttmästaren
och
Riddaren
Hildebrand
,
varit
sinnad
,
att
låta
dagsverkare
vid
kyrkotakets
täckande
få
en
liten
dagspeng
ur
kyrkans
kassa
;
men
vid
närmare
övervägande
har
Högbem:te
Patron
funnit
kassan
så
svag
,
att
den
icke
mäktar
bestrida
utgifterna
för
Spån
och
Spik
och
avbetalningen
till
Byggmästaren
.

Såsom
ock
församl
:
n
varnades
,
att
hysa
och
giva
något
åt
de
så
kallade
häktmakare
och
dylika
.
§
31
.

Lind
,
att
benäget
besörja
om
dessa
järnplåtars
förfärdigande
och
om
oljans
förskaffande
;
vilket
lovades
.
2:o
.

Sockenmännen
Pär
i
Harstorp
betalade
nu
sin
skuld
med
räntan
till
kyrkokassan
.

Församl
:
n
beslöt
,
att
gl.
Pigan
Kerstin
i
Tyblenäs
skulle
få
intaga
det
lediga
rummet
i
fattgstugan
.
§
8
.

Lind
trodde
,
det
hans
Herre
icke
heller
skulle
vara
däremot
.

Uppläst
och
till
alla
delar
vidkänt
,
betyga
Johan
Lind
P
.
Diuhlstedt
Peter
Petersson
i
Brenäs
Jonas
Jonsson
i
Trolldal
nämndeman
Bängt
Pärsson
i
Remröd
Sexmän
År
1785
den
8
Maj
,
efter
vanlig
pålysning
,
blev
allmän
Valborgsmässo
Sockenstämma
hållen
med
St.
Malms
församl
.
,
i
närvaro
av
vanliga
Herrskapens
Betjänter
och
Sockenmän
,
på
följande
vis
:
§
1
.

Till
takfotens
bestrykande
på
kyrkan
i
sommar
föreslog
klockaren
och
målaren
Nyhlin
,
utom
det
förråd
kyrkan
därav
äger
förut
,
ännu
3
kannor
olja
och
IV2
pund
blivit
,
varvid
församl:s
Invånare
erinrade
,
att
då
skulle
även
muras
under
fjärbräderna
på
västra
gaveln
.
§
4
.

Föregående
2:ne
Protokoll
erkännas
till
alla
delar
betyga
Gerhard
Lind
P
.
Djuhlstedt
Erik
Andersson
i
Mogetorp
Jonas
Olsson
i
Walla
Sexmän
Peter
Petersson
i
Brenäs
nämndeman
År
1786
d
.
25
Maj
,
efter
förut
skedd
tillräcklig
pålysning
,
blev
ordentl.
Valborgsmässo
Sockenstämma
med
St.
Malms
församl
.
hållen
,
i
närvaro
,
å
välborne
Herr
Patroni
vägnar
,
av
Bruksinspektorn
Herr
Gerhard
Lind
,
å
St.
Djulö
respektive
ägare
,
av
frälse
Befall
.

Församlingen
anmodade
Sexman
i
Valla
,
att
detta
arbete
om
måndag
sig
åtaga
och
begynna
,
vilket
lovades
,
och
Sexman
i
Stensjö
fick
tillsägelse
att
därtill
bestyra
om
sprängd
stens
framskaffande
,
som
fanns
vid
Brogtorp
.
§
5
.

Pastor
varnade
alla
dem
,
som
komma
att
gräva
åt
lik
,
att
de
icke
skola
låta
de
dödas
ben
ligga
ovan
jord
,
som
kunna
bli
uppkastade
vid
grävningen
,
utan
,
så
snart
ett
lik
är
nedsatt
och
jordfäst
,
böra
de
först
nedkasta
de
uppgrävna
ben
och
huvudskallar
och
sedan
mullen
därpå
.
§
7
.

Vid
sista
Prästmötet
avgjordes
,
att
när
kommunion
hålls
i
en
kyrka
,
så
skall
hela
församl
:
n
stå
uppe
,
medan
kommunion
påstår
,
och
kyrkodörrarna
skola
igenstängas
,
när
syndabekännelsen
läses
och
de
allmänna
skriftermålen
hållas
,
på
det
deras
andakt
,
som
inne
är
,
ej
må
störas
av
de
inkommandes
buller
.
:
vilket
Pastor
nu
kungorde
till
allas
efterrättelse
.
§
12
.

Ingen
var
,
som
icke
härtil
gav
sitt
samtycke
och
bifall
,
utlovandes
att
det
efterkomma
.
§
15
.

Men
som
2
Sexmän
är
på
Djula
gods
,
vilka
äga
dagsverksfrihet
,
ty
av
gå
3A
mantal
,
resten
således
193
/
s
och
dagsverken
högst
19
för
jämn
räkning
må
det
dock
förbli
vid
20
dagsverken
uti
vart
skov
och
täcktes
herr
kyrkoherden
och
församling
varje
söndag
tillsäga
Sexm.
Jonas
i
Trolldahl
,
vilka
dagar
Djula
gods
bör
sig
infinna
i
Prästagn
.

Lind
,
Pastor
tillsporde
Sexmännen
,
varför
de
icke
ville
göra
dagsverken
vid
prästgårds
Byggnaden
,
sedan
de
flera
resor
blivit
tillsagda
därom
,
helst
ingen
förordning
befriar
dem
därifrån
?

Maj:t
allernådigast
dem
erbjudna
husbehovsbränningen
?

Maj:ts
nådiga
befallning
utfärdade
Kungörelser
,
angående
en
fri
husbehovsbrännings
arrenderande
av
Socknens
Invånare
,
får
jag
härmed
förklara
det
jag
för
de
av
mig
i
Socknen
ägande
Säterier
,
med
därtill
lydande
rå-
och
rörscheman
,
så
väl
som
de
hemman
,
vilka
jag
har
under
noga
bruk
,
alldeles
avsäger
mig
samma
i
nåder
erbjudna
arrende
,
och
vad
mina
i
Socknen
belägna
frälsehemman
som
av
bönder
brukas
,
angår
,
så
må
det
ankomma
på
åbornas
eget
fria
val
att
därutinnan
göra
,
som
de
för
sig
bäst
och
nyttigast
finna
;
dock
med
det
kraftiga
förbehåll
å
min
sida
,
att
vad
de
härutinnan
göra
eller
låta
,
aldrig
annorl
.
må
anses
än
såsom
en
deras
egen
personl
.
förbindelse
som
med
mina
hemman
ingen
gemenskap
äger
,
och
för
vars
uppfyllande
samma
hemman
varken
nu
eller
i
tillkommande
tider
kunna
häfta
;
ävensom
jag
ock
förbehåller
mig
att
hos
åborna
och
uti
dess
egendom
njuta
den
förmånsrätt
för
innestående
avrad
och
husröteandel
,
som
allmänna
lagen
jordägare
och
räntegivare
tillägger
,
i
fall
åbon
eller
skattebonden
skulle
brista
i
det
kontrakt
han
med
Kungl.
Maj:t
och
Kronan
ingår
.

Därefter
tillspordes
skattebönderna
,
vad
beslut
de
fattat
i
förevarande
ämne
?

Efter
uppläsandet
härav
begärde
Befallningsmannen
Djulstedt
del
av
denna
uträknig
,
för
att
kommunicera
den
med
Kammarherren
välborne
Herr
C
.
Uggla
;
vilket
bifölls
,
med
åstundan
,
att
få
Hr
Kammarherrens
svar
härpå
nästa
söndag
.

År
1787
d
.
4
Nov
.
inkallades
Socknens
Invånare
i
Sockenstugan
,
då
Pastor
frågade
,
om
någon
vore
närvarande
från
Djula
,
att
avgiva
svar
,
angående
den
i
dag
8
dar
sedan
uppläst
uträkningar
om
fönster
i
Prästgården
?

Nu
beslöts
således
,
att
vart
matlag
skall
i
stället
för
6
giva
8
runstycken
.

Alm
och
hans
hustru
framkom
och
berättade
,
att
så
snart
de
fann
sin
son
död
,
har
de
budat
till
sig
Bonden
Pehr
Pehrsson
och
änkan
Kerstin
Simonsd:r
i
Kårtorp
,
vilka
strax
inställde
sig
.

Som
församlingens
Patronus
,
Ryttmästaren
och
Riddaren
välborne
Hr
David
Hildebrand
bifallit
detta
byte
utan
något
förbehåll
,
men
Kammarherren
välb.
Herr
Carl
Uggla
samtyckt
därtill
med
villkor
,
att
samma
hus
skulle
säljas
på
auktion
;
så
frågade
Pastor
,
om
församlingens
vilja
vore
att
de
skulle
auktioneras
och
varpå
svarades
:
ja
.

Boken
måtte
intagas
så
lydande
:

Till
övre
Våningen
:
9
tolfter
plank
till
golv
ven
å
24
d:r
12
Dito
bräder
till
panel
å
14
d:r
6
dörrkarmar
å
9
d:r
6
dörrar
å
18
d:r
13
St.
fönsterkarmar
å
12
d:r
52
St.
fönsterbågar
å
IV2
d:r
52
St.
fönster
fotpanelning
i
5
rum
å
12
d:r
6
par
dörrgångjärn
å
3
d:r
beslag
till
13
fönsterluckor
å
14
d:r
6
st.
polerade
dörrlås
å
9
d:r
5
Segelgarn
till
gipsningen
å
3
d:r
18
tjog
oskalad
rönn
till
taken
å
6
d:r
13250
St.
gipsspik
å
9
d:r
Rummens
vitlimning
med
kosthållning
Snickare
arbetat
med
golv
etc.
5
St.
gröna
Kakelugnar
med
uppsättning
å
84
d:r
hemförseln
från
Nyköping
Kakelugnsmakares
kost
under
uppsättningen
5
St.
dubbla
Kakelugnsdörrar
å
24
d:r
5
St.
Kakelugnsfötter
å
20
d:r
5
St.
gjutna
Spjäll
å
9
d:r
13
St.
vattenbläck
till
fönsterna
5
St.
Kakelugnspipor
av
plåtar
Målaren
för
dörrar
och
dörrfoders
med
fönsterkarmars
och
bågars
samt
vattenbläckens
överstrykning
med
oljefärg
,
efter
räkning
Till
nedre
våningen
:
12
—
9
16
.
3
—
6
—
8
32
.
4
16
.
42
40
.
3
16
.
1
—
10
5
.
4
.
3
—
40
.
6
—
6
.30
.
1
:
32
.
8
:
14
.
8
.
23:16
.
2:24
.
1:43
.
6:32
.
5:26
.
2:24
.
2:16
.
—
:
45
.
7
:
—
.
6
St.
Ekbjälkar
till
dörrkarmar
i
förstugan
2:24
.
2
St.
gröna
Kakelugnar
å
84
d:r
9:16
.
dessas
transport
från
Nyköping
—
40
.

Pehr
i
Smedstorp
anmälde
vidare
,
att
drängens
tokiga
moder
,
som
sitter
i
hus
därstädes
,
skall
mycket
vara
orsaken
till
Sonens
täta
besök
i
Smedstorp
,
helst
hon
går
in
till
hospitalet
och
lockar
honom
ut
med
sig
.

Med
överläggning
av
detta
ämnet
uppsköt
församlingen
till
en
annan
gång
.
6:o
Beslöts
,
att
gamla
Sockenstugetimret
skulle
nu
i
veckan
sönderhuggas
åt
de
fattiga
till
ved
av
dem
,
som
annars
vore
i
ordning
,
att
till
fattighuset
framskaffa
ved
.
7:o
Bifölls
,
att
till
eldning
i
Sockenstugan
om
Söndagsmorgnarna
vintertiden
böra
årligen
3
å
4
lass
huggen
ved
framköras
på
samma
sätt
,
som
i
föregående
6
§
nämnt
är
.
8:o
Avgjordes
att
Kyrkbacken
skulle
med
första
öres
)
av
alla
8
rotarne
,
några
var
dag
,
tills
den
blev
fullärd
.
9:o
Nämndemännen
anmodades
,
att
utlysa
och
hålla
auktion
på
gamla
fönster
,
järn
och
spik
,
som
suttit
i
gl.
Sockenstugan
.
10:o
De
resterande
med
fattigdelen
för
1788
uppnämndes
och
tillsades
,
att
den
ofördröjligen
betala
.

De
förmanades
,
att
härpå
ha
noga
akt
,
på
det
att
ordning
och
skick
i
Guds
hus
må
bibehållas
.

Maj
1790
uppläste
,
och
riktigheten
därav
erkänt
betyga
Gerhard
Lind
A
.
Blomberg
Pehr
Pehrsson
i
Brenäs
nämndeman
Olof
Pärson
i
Banninge
Eric
Andersson
i
Walla
Kyrkovärdar
Jonas
Erickson
i
Walla
Erick
Pärson
i
Remröd
Sexmän
År
1790
d
.
9
Maj
,
efter
14
dagars
förut
skedd
pålysning
,
blev
allmän
Valborgsmässo
Sockenstämma
med
St.
Malms
församl
.
hållen
,
i
närvaro
av
resp
.

Lind
ingav
till
Malms
församl
.
för
Socken
och
fattigstugebyggnaden
en
räkning
på
302
R
.
36
s.
11
rst
.
,
som
upplästes
och
erkändes
.

Kajsa
Pehrsd:r
i
Heden
blev
intagna
i
3:dje
fattigklassen
,
samt
Pig.
Maja
Simonsd:r
i
Kärtorp
uti
den
2:dra
klassen
.

Lind
i
sista
Sockenstämman
givit
,
angående
Magasins
husets
försäljande
till
hjälp
vid
betalningen
för
Socken
och
fattigstugebyggnaden
,
gav
bem:te
H:r
Inspektor
strax
vid
handen
,
att
S
.
T.19
)
herr
Patronus
för
sin
del
bifaller
Magasinshusets
försäljande
.

Juli
1789
gjorde
och
efter
bemälda
Befallningsmans
död
hos
Oppunda
Häradrätts
vid
förlidna
)
års
höstting
den
)
27
Nov
.
(
ember
)
1794
behörigen
vigilerade
Testamente
updragit
mig
en
oinskränkt
rätt
samt
fullmakt
och
myndighet
,
att
om
dess
efterlämnade
kvarlåtenskap
disponera
och
giva
densamma
,
antingen
hel
och
hållen
eller
delad
,
åt
vem
eller
vilka
mig
skulle
nyttigast
synas
,
samt
jag
till
följa
därav
föranstalta
låtit
,
dels
att
den
avlidnes
mindre
betydliga
kvarlåtenskap
av
Kläder
och
annat
kommit
till
något
gagn
åt
hans
mest
älskade
vänner
och
sådana
i
behov
varande
,
som
närmast
stått
under
hans
lydnad
och
honom
till
nöjes
samt
med
tillgivenhet
sig
uppfört
,
dels
att
hans
redbarare
egendom
blivit
efter
dess
högsta
möjliga
värde
förvandlad
,
varvid
densamma
jämte
de
i
hans
Bo
befintliga
kontanta
penningar
tillsammans
utgjort
en
summa
,
vilken
då
därtill
läggas
så
väl
den
ränta
jag
därpå
kunnat
uppbringa
till
den
lista
i
denna
månad
,
som
något
mera
,
vartill
,
att
dessa
medel
föröka
,
utvägar
under
den
förflutna
tiden
för
mig
sig
yppat
,
bestiger
sig
i
Riksgäldssedlar
till
ett
Kapital
stort
Ett
Tusende
fem
Hundrade
Trettio
Tre
Riksdaler
Sexton
skilling
/
:
1533
Rdr
16
s
:
/
;
så
har
jag
vid
mitt
fattade
beslut
om
dessa
pgrs
(
penningars
)
användande
med
desto
större
nöje
och
tillfredsställelse
funnit
mig
både
skyldig
och
villig
att
giva
uppmärksamhet
åt
Testatorns
i
livstiden
oftast
för
mig
muntligen
i
denna
delen
yttrade
åstundan
,
som
därigenom
vardar
ett
välgörande
och
honom
hedrande
kristendomsverk
befordrat
;
och
förordnar
jag
fördenskull
härmedelst
,
att
av
ovannämnde
Kapital
1533
Rdr
16
s
(
sk
)
riksgälds
Sedlar
skola
.
lo
Tre
Hundrade
Trettio
Tre
Riksdaler
16
s
(
sk
)
/
:
333
R
.
16
:
/
Riksgälds
sedlar
med
6
procents
ränta
därpå
från
den
1
sta
nästlidne
)
Maj
till
samma
tid
nästa
år
1796
då
överlämnas
till
Lasarettet
i
Nyköpings
Stad
,
att
jämte
de
övriga
Lasarettsmedlen
användas
till
där
inkommande
sjuklingars
underhåll
,
läkemedel
och
hjälpsammaste
omvårdnad
;
varvid
med
den
säkra
förmodan
jag
hyser
att
dessa
angivna
medel
under
Lasaretts
Direktionens
ömma
och
sorgfälliga
omsorg
på
bästa
sätt
i
sitt
ändamål
disponeras
och
användas
,
jag
blott
gör
det
förbehåll
,
som
själva
erkänslan
för
denna
undfångna
gåvan
villigen
och
genast
lär
rättfärdiga
,
att
nämligen
en
billig
företrädes
rätt
lämnas
dem
från
Ericsbergs
gård
med
tillydande
Hemman
och
lägenheter
,
vilka
under
den
tid
min
Käre
)
Son
,
välborne
)
Herr
David
Gotthard
Hildebrand
denne
egendom
innehar
,
kunna
komma
i
den
ömkansvärda
belägenhet
,
att
vara
nödsakade
inom
Lasarettet
söka
räddning
för
sitt
liv
och
hälsa
.
2o
de
övriga
Ett
Tusende
Två
Hundrade
/
:
1200
:
/
Riksdaler
Riksgäldssedlar
vara
med
nedannnämnda
villkor
och
under
förbehåll
,
att
de
noga
efterlevas
,
givna
till
St.
Malms
Församlings
fattig
Kassa
och
skola
under
bemälde
min
K
.
(
är
)
Sons
Herr
David
Gotthard
Hildebrands
livstid
bli
hos
Honom
innestående
emot
Sex
procents
ränta
,
men
när
min
K
.
(
är
)
Son
död
är
,
bör
det
som
av
ovanberörda
Kapital
1200
Rdr
kan
vara
övrigt
,
genast
avlämnas
till
St.
Malms
församlings
fattig
Kassas
Föreståndare
,
vilka
med
laga
ansvar
och
i
samråd
med
Possessoren
av
Ericsbergs
fidei
commiss
äga
att
besörja
,
det
,
de
då
undfängna
medlen
vara
med
största
möjliga
)
säkerhet
och
till
bästa
förmån
förräntade
,
samt
för
övrigt
då
vaka
även
därpå
,
att
berörda
gåva
rätteligen
efter
detta
förordnande
användas
.
—
Som
Ericsbergs
gods
underhavande
inom
St.
Malms
Socken
och
bland
dem
i
synnerhet
den
torftigare
delen
,
under
Testators
uti
berörda
Socken
in
till
dess
död
tillbringade
mångåriga
levnad
,
alltid
ägt
förnämsta
föremålet
för
dess
ömhet
och
omvårdnad
,
så
bör
efter
dess
önskan
,
den
jag
jämväl
härutinnan
gärna
efterföljer
,
varken
nu
eller
framledes
några
andra
kunna
komma
att
njuta
understöd
och
hjälp
av
ovannämnde
förlänta
och
donerade
medel
,
eller
därav
få
sig
begagna
,
än
sådana
gamla
,
orkeslösa
,
fattiga
och
sjukliga
,
jämte
värnlösa
barn
,
vilka
eller
vilkas
föräldrar
längre
tid
tjänat
och
arbetat
under
Ericsbergs
gods
,
samt
är
på
de
under
Ericsbergs
gård
inom
St.
Malms
Socken
lydande
hemman
och
ägor
boende
,
samt
under
föregående
levnaden
gjort
sig
kända
för
gudsfruktan
,
redligt
och
beskedligt
uppförande
samt
arbetsamhet
;
och
då
antalet
av
dylika
nödställda
icke
bör
bli
stort
,
därest
efter
min
hägnesamma
förhoppning
Ericsbergs
Possessoren
framledes
och
i
den
påföljande
tiden
såsom
nu
med
efterföljd
av
det
lovvärda
efterdöme
den
avlidne
Instiftaren
av
Ericsbergs
fideicommiss
under
sin
levnad
givit
,
låter
sig
ömmast
om
hjärtat
ligga
,
att
mot
sitt
folk
vara
en
öm
Fader
och
välgörande
husbonde
,
som
gärna
av
sitt
eget
förråd
efter
omständigheterna
hjälper
en
i
nöd
och
behov
kommen
trogen
,
redlig
och
flitig
tjänare
,
finner
jag
både
för
gott
och
lämpligast
,
att
antalet
av
dem
,
vilka
efter
denna
2
§
i
detta
mitt
förordnande
och
av
där
givna
Kapitalet
komma
att
njuta
underhåll
,
bör
inskränkas
inom
Tio
/
:
10
:
/
till
högst
Femton
/
:
15
:
/
de
mest
behövande
,
vilkas
utnämnande
,
jämlikt
de
grunder
jag
nu
utstakat
,
helt
och
hållet
ensamt
och
ovillkorligen
skall
ankomma
nu
och
framledes
på
Ericsbergs
Possessors
gottsinnande
och
val
,
efter
de
behövliga
underrättelser
han
så
väl
av
Pastor
i
St.
Malms
församling
)
som
andra
vederbörande
var
till
sin
upplysning
inhämtande
;
såsom
jag
ock
Ericsbergs
Possessor
gemensamt
med
Pastor
i
St.
Malms
(
församling
)
och
denna
Sockens
fattigkassas
föreståndare
uppdrager
och
förbinder
,
att
med
all
oförtrutan
omsorg
vaka
och
tillse
,
det
understödet
till
det
belopp
,
som
här
nedanför
stadgas
,
årligen
,
så
länge
något
av
det
givna
Kapitalet
är
övrigt
,
riktigt
utgår
och
kommer
till
hända
åt
de
personer
,
vilka
årligen
utnämnas
att
bli
delaktiga
av
samma
understöd
,
däruti
de
undfå
vardera
en
efter
vars
och
ens
omständigheter
,
nöd
och
belägenhet
,
som
Ericsbergs
Possessor
ensamt
äger
att
pröva
,
proportionerad
andel
,
som
dock
för
någon
må
ej
överstiga
eller
bli
större
än
en
Femte
del
/
iVs
:
/
och
icke
eller
för
någon
bli
mindre
än
en
Tjugondel
/
:

Inlämnades
och
upplästes
följande
Räkning
:

Jonas
i
Heden
yrkade
åter
,
å
grannens
smedens
och
dess
hustrus
i
Heden
vägnar
,
som
för
ålderdoms
bräckligheter
i
dag
ej
kunde
vara
närvarande
,
att
de
måtte
i
fattighuset
intagas
.

Församlingens
beslut
blev
,
att
de
skulle
få
2
skilling
)
för
paret
av
de
personers
skor
,
som
är
äldre
och
mantalsskrivna
,
men
1
skilling
)
6
runstycken
för
paret
av
de
personers
skor
,
som
är
yngre
och
ej
kommit
i
mantal
.
§
8
.

Men
den
4des
man
yttrade
sig
kunna
förse
sin
hustru
med
nödigt
uppehälle
.
§
4
.

Eric
Nilsson
i
Prästorp
och
Jan
Olsson
i
Horssnäs
antogs
till
sexmän
,
den
förre
i
Kyrko
och
den
senare
i
Bålsnäsrotar
,
uti
deras
ställe
,
som
begärt
avsked
.
§
6
.

Både
han
och
sådana
kreaturs
ägare
undfick
nu
eftertryckl
.
(
iga
)
föreställningar
,
att
lagen
i
detta
mål
noga
åtlyda
.

Under
anmälan
,
det
skall
allmogen
i
nästgränsande
socknar
ha
vid
hållna
sockenstämmor
överenskommit
,
att
hos
Konungens
Befallningshavande
i
länet
anhålla
,
det
ville
Konungens
Befalln
.
(
ingshavande
,
i
anseende
till
svårigheten
och
kostnaden
för
allmogen
vid
sina
soldaters
utrustande
till
regementsmöten
,
hos
Kgl.
Majestät
underdånigast
hemställa
,
det
kunde
för
i
år
,
då
sådan
dyrhet
är
å
både
ätande
och
tärande
varor
,
allmogen
i
nåder
lisas
från
)
det
regementsmöte
,
vilket
,
efter
vad
de
hört
,
skulle
fram
på
sommaren
komma
att
hållas
med
Söderm
.
(
anlands
)
Kgl.
infanteriregemente
;
har
en
del
av
St.
Malms
sockenbor
av
allmogen
begärt
,
det
måtte
församl
.
(
ingens
invånare
inkallas
i
sockenstugan
,
för
att
i
enahanda
ämne
få
samrådas
.

Välborne
Herr
Patronus
täcktes
själv
tillkännagiva
,
att
genom
ett
utav
avl
.
(
idne
)
Brucks
Inspektorn
Taxels
Änka
,
Anna
Maria
Vinter
,
vid
Cathrineholm
,
gjort
Testamente
av
d
.
(
en
)
6
.

Slutligen
)
beslöts
,
det
sockenstämmo
protokoll
häröver
skulle
upprättas
,
för
att
till
K
.
(
ungliga
)
patriotiska
sällskapet
insändas
tillika
med
det
skriftl
.
(
iga
)
betyget
.

Okt
.
(
ober
)
hölls
allmän
Mickelsmässo
Sockenstämma
med
St.
Malms
resp
.
(
ektive
)
församl
.
(
ing
)
.
§
1
.

Efter
noga
undersökning
,
varav
det
härrörde
,
att
det
inre
i
klockstapeln
var
sviktande
under
ringningarna
,
befanns
det
komma
därav
,
att
viggarna
under
bjälkarne
var
multnade
och
inre
muren
,
varpå
underslaget
vilar
,
något
sjunken
.

Notarien
i
Kgl.
Svea
Hovrätt
Herr
Anders
Lindblad
och
kyrkov
.
(
ärden
)
i
Stensiö
Pehr
Ersson
utsedde
och
förordnade
,
att
i
detta
mål
vara
socknens
ombud
och
dess
rätt
och
bästa
bevaka
.

Oktober
blev
efter
ordentlig
)
pålysning
,
i
närvaro
av
församlingens
Herr
Patronus
och
Sockenmännen
,
den
allm
.
(
änna
)
Mickelsm
.
(
ässo
)
Sockenstämma
med
St.
Malms
församling
)
hållen
.
§
1
.

Särskilt
stolrum
i
Kyrkan
ville
man
tills
vidare
ej
bevilja
sockenhantverkare
,
utan
må
de
sitta
i
deras
bänkar
,
vars
hushjon
de
är
,
eller
söka
sig
rum
i
de
nya
bänkarna
.
§
8
.

Förlidet
år
hade
Ridder
åter
utan
församlingens
lov
med
sina
anhöriga
inkommit
i
församl
.
(
ingen
)
och
satte
sig
i
hus
på
förr
nämnda
ställe
,
varom
undertecknad
genom
upplästa
skrivelsen
fick
kunskap
,
som
befallde
sexman
av
visa
denna
Ridder
ur
församl
.
(
ingen
)
varå
Ridder
skall
gyckelaktigt
svarat
,
att
han
väl
skulle
begiva
sig
bort
,
allenast
undertecknad
kunde
skaffa
honom
något
bättre
,
då
han
ville
färdas
och
taga
stugan
med
sig
.

Och
som
förmärktes
,
att
större
delen
av
dessa
uppnämnde
fattiga
och
i
de
frånvarandes
ställe
deras
närmaste
anhöriga
var
nu
tillstädes
;
så
tillsades
,
att
om
de
ville
dröja
kvar
,
till
dess
sockenstämman
blivit
slutad
,
så
skulle
de
i
dag
undfå
hälften
av
den
dem
beviljade
pgr
summa
,
men
den
andra
hälften
ej
förr
än
vid
Olofsmässan
)
;
hkt
(
vilket
)
ock
skedde
.
§
3
.

Listan
på
de
15
fattiga
,
som
respektive
Possessorn
av
Ericsberg
för
i
år
behagat
utnämna
till
åtnjutande
av
100
Rdr
,
upplästes
.
§
4
.

Sexman
i
Löpsjötorp
frågade
,
om
sängliggande
hustrun
i
Charlottendal
kunde
ur
fattigkassan
få
pgr
.
(
penningar
)
till
läkemedel
för
sin
sjukdom
?

Emellertid
fick
de
allvarliga
)
tillsägelser
,
att
icke
besvära
någon
socken
utom
Malm
med
tiggande
.
§
6
.

Änk
.
(
an
)
Kerstin
Månsdotter
i
Korsshellstugan
)
och
flickan
Ulla
Pehrsdotter
i
Löskbol
anmäldes
såsom
de
där
ärna
i
sommar
dricka
Medevi
brunn
,
med
begäran
om
fattigdoms
bevis
.

In
fidem
C
.
F
.
Maneck
Uppläst
och
erkänt
:

Landshövdingens
fullmakt
.
§
7
.

Och
så
snart
hon
då
märkte
barnet
vara
dött
,
bad
hon
sin
man
inkalla
först
änkan
Stina
Håkansdotter
och
sedan
hustrun
Anna
Maja
Taberman
vid
Forssjö
,
att
upptaga
och
bese
barnet
.

I
dag
fick
ur
fattigkassan
följande
torftiga
personer
pgr
.
(
penningar
)
:

Sockenmännen
stannade
i
det
beslut
,
att
Klingström
skulle
befrias
från
böter
och
magen
,
om
nämndeman
ville
antaga
honom
till
dräng
,
få
vara
i
församlingen
.

Enligt
förlidet
års
beslut
skulle
emellertid
taken
över
bodar
och
brygghus
i
Prästgården
nästa
vecka
med
torv
och
näver
repareras
,
även
som
skulle
över
stallet
då
förbättras
med
2
polster
sågbakar
för
32
s
(
sk
)
Banco
,
vartill
kyrkokassan
för
församlingen
skulle
gå
i
förskott
.
§
10
.

Sockenmännen
varnades
,
att
icke
bortslösa
sin
spannmål
genom
överflödigt
brännvinsbrännande
och
supande
.
§
8
.

Lars
Nilsson
,
såsom
sexman
i
den
roten
,
ålades
,
att
ännu
en
gång
allvarligen
påminna
Pehr
Andersson
att
förfoga
sig
ur
socknen
,
och
i
händelse
Pehr
Andersson
ej
efterkommer
denna
slutliga
varning
,
skulle
man
omsider
genom
kronobetjäningen
vidtaga
tjänliga
mått
och
steg
.
§
7
.

Räkningen
uppgick
,
tegel
,
kalk
,
plank
,
bräder
,
spik
,
järn
oberäknat
,
till
ett
belopp
i
penningar
av
femtio
fem
Riksdaler
,
47
skill
.

Riksgäldsmynt
,
vilka
Herr
Friherre
Bonde
på
Ericsberg
för
församlingen
utgivit
,
och
komma
att
,
sammanlagda
med
vad
den
ännu
ouppgjorda
räkningen
för
tegel
,
kalk
,
plank
,
bräder
,
spik
,
järn
,
som
även
bemälde
Herre
till
reparationen
för
församlingen
lämnat
,
innehåller
,
till
betalning
på
församlingen
lämnat
,
innehåller
,
till
betalning
på
församlingen
reparteras
.

Den
ovannämnde
räkningen
tillika
med
kvittenserna
och
penningar
beloppet
55
Riksdaler
,
47
skil
.

Riksgäldsmynt
godkändes
till
alla
delar
av
Församlingen
.

Sålunda
vara
avgjort
och
beslutat
;
intyga
å
församlingens
vägnar
undertecknade
:

E
.
Folien
kyrkoherde
År
1812
den
6te
december
ankom
till
kyrkan
och
upplästes
från
predikstolen
Höglovlige
)
Lands
Hövdinge
Ämbetets
kungörelse
om
skatt
skrivningen
med
St.
Malms
Socken
den
21
och
22
December
1812
,
då
även
Kungl
.

Majts
Förordning
av
den
30
September
1812
angående
mantals
och
skattskrivningarna
i
Riket
från
predikstolen
upplästes
,
varjämte
församlingen
inlystes
i
sockenstugan
,
varest
Landshövdinga
Ämbetets
ovansagde
kungörelse
för
församlingen
omlästes
.

Och
sedan
Anno
etc.
72
under
salig
Konung
IAHANS
Regering
,
i
Upsala
allmänna
Prästmöte
på
nytt
bekräftat
.

Sonen
är
av
Fadern
allena
,
icke
gjord
,
icke
skapat
,
utan
född
.

En
är
han
,
dock
icke
så
,
att
Gudomen
är
förvandlat
i
mandomen
,
utan
Gudomen
har
till
sig
annamat
mandomen
.

Var
ock
det
ordet
PERSON
,
hos
oss
brukat
uti
samma
märkelse
,
som
de
gamla
Församlingarnas
Lärare
,
i
denna
saken
det
brukat
har
,
Nämligen
,
att
det
märker
icke
någon
del
eller
egenskap
uti
andra
;
utan
det
som
egentligen
är
och
sin
varelse
har
i
sig
själv
.

Item
,
de
Valentinianer
,
Arrianer
,
Eunomianer
,
Mahometister
och
andra
slika
.

Den
samma
Christus
skall
ock
uppenbarligen
komma
,
till
att
döma
levande
och
döda
,
etc.
efter
den
Apostoliska
Tros
Bekännelsen
.

ATT
vi
denna
Tro
måtte
bekomma
,
är
Predikoämbetet
instiftat
,
genom
vilket
Evangelium
förkunnas
,
och
Sakramenten
utdelas
.

Ifrån
de
fördolda
synder
rena
mig
.

De
vara
ock
så
undervisade
,
att
alla
människostadgar
,
som
är
instiftade
till
att
blidka
Gud
,
förtjäna
Guds
nåder
,
och
tillfyllestgöra
eller
betala
för
synderna
,
är
tvärt
emot
det
helga
Evangelium
,
och
Trons
lära
.

Och
skall
hela
denna
läran
om
Tron
,
bli
brukat
emot
den
strid
och
kamp
,
som
förskräckt
samvete
plägar
vederfaras
,
och
utan
sådana
samvets
kamp
kan
hon
intet
rätt
bli
förstånden
.

Och
Guds
Församling
sjunger
:

Allenast
bortlägger
de
några
missbruk
,
vilka
är
nya
,
och
emot
den
grund
och
mening
,
som
Canones
,
eller
den
gamla
Kyrkolagen
innehåller
,
av
olärde
och
onde
lärare
upptagna
:

Själve
Canones
eller
Kyrko
lagen
,
medgiver
ock
,
att
man
väl
må
understundom
uti
efterkommande
tider
för
mänsklig
svaghet
skull
,
lindra
den
gamla
strängheten
.

Sammaledes
råder
ock
Cyprianus
,
att
de
kvinnor
som
icke
hålla
kunna
den
utlovade
kyskheten
,
må
giva
sig
i
mans
våld
.

Desslikes
behålles
ock
något
så
när
alla
brukliga
Ceremonier
,
allenast
att
ibland
Latinska
Sånger
var
somligstädes
Sånger
på
eget
tungomål
brukade
,
vilka
tillagda
är
,
folket
till
att
lära
och
undervisa
.

Folket
blir
ock
tillvant
,
att
de
ock
tillika
gå
till
Herrens
Nattvard
,
om
några
där
ibland
är
skickliga
:
vilket
ock
förökar
Religionen
,
och
vyrdningen
emot
de
allmänneliga
Ceremonier
och
stadgar
.

Där
till
med
som
ock
den
mening
,
som
har
så
förökat
hemliga
Vråmässor
,
att
de
är
otaliga
vordna
,
nämligen
,
att
Christus
med
sitt
lidande
har
fyllestgjort
och
betalt
för
Arvssynden
,
och
sedan
förordnat
Mässan
,
uti
vilka
skulle
ske
offer
,
för
dagliga
synder
,
så
väl
grova
,
som
de
av
svaghet
hända
är
.

Där
till
med
,
uppläses
den
helga
Skrift
,
uti
den
Staden
Alexandria
,
var
Onsdag
och
Fredag
,
och
de
förnämligaste
Lärare
har
henne
uttytt
,
och
all
ting
förhandlat
där
förutan
någon
Mässa
.

Ty
det
är
många
synder
som
man
varken
förstå
eller
minnas
kan
.

Till
det
första
,
är
den
läran
om
Guds
nåd
och
den
rättfärdighet
som
kommer
igenom
Tron
,
mycket
förmörkat
,
vilken
är
den
förnämste
del
av
Evangeliet
,
och
bör
alltsommest
driven
och
predikat
bli
i
Guds
Församling
,
på
det
att
Christi
förskyllan
måtte
alla
väl
kunnig
vara
,
och
Tron
som
tror
synderna
förlåtas
för
Christi
skull
,
kunna
långt
över
gärningarna
räknat
bli
.

Och
man
har
menat
,
att
hela
Kristendomen
skulle
stå
där
uti
,
att
man
höll
vissa
Helgdagar
,
vissa
Stadgar
,
Fastedagar
och
Klädbonad
.

De
indraga
ock
vittnesbörd
av
den
helga
Skrift
:

Item
,
Efter
ni
nu
döda
är
med
CHristo
,
ifrån
de
världsliga
stadgar
,
vi
låter
ni
er
då
begripas
med
beskrivna
stadgar
?
lika
som
ni
ännu
lever
i
världen
,
de
där
säga
,
du
skall
icke
komma
vid
det
,
icke
smaka
det
,
icke
hantera
det
.

Här
förkastar
våra
motståndare
oss
,
att
våra
Lärare
förbjuder
köttets
tvång
och
aga
,
vilket
den
Kättaren
Iovianus
i
förtiden
lärt
har
.

Åtskillnad
på
Fastedagar
syndrar
icke
Trons
enighet
:

Vad
om
Klosterlöften
hos
oss
lärt
var
,
kunna
de
samma
bättre
befinna
och
förstå
,
som
minnas
vad
skick
uti
Klostren
varit
har
,
och
hur
mycket
där
inne
dagligen
är
gjort
och
bedrivit
emot
den
gamla
Kyrkolagen
.

Till
dessa
villfarelser
har
och
kommit
en
sådan
mening
om
Klosterlöften
,
den
ock
i
förtiden
själva
Munken
,
som
något
förståndigare
vore
,
misshagat
har
:

Det
kan
icke
heller
nekas
,
att
Munkarna
har
ju
lärt
,
sig
genom
Klosterlöften
och
andra
sådana
sina
stadgar
bli
rättfärdiga
,
och
förtjäna
syndernas
förlåtelse
,
Ja
,
de
har
uppdiktat
grovare
villfarelser
,
i
det
de
säga
sig
kunna
meddela
andra
sina
gärningar
.

Dessförinnan
i
utvärtes
måtto
flitigt
göra
goda
gärningar
,
och
akta
sitt
stånd
och
ämbete
.

Om
sådana
saker
är
mycket
av
nöden
förmana
folket
.

Ty
det
andliga
Regementet
har
sina
synnerliga
befallning
till
att
predika
Evangelium
och
utskifta
Sakramenten
.

De
införa
ock
Apostlarnas
exempel
uti
Apostla
Gärningarna
,
i
det
15
Kap:
Där
de
har
förbjudit
äta
blod
,
och
det
som
var
förkvavt
.

Men
det
är
uppenbart
,
att
människo
stadgar
är
för
sådana
falsk
mening
skull
,
otaliga
många
vordna
i
Församlingarna
,
och
den
läran
som
är
om
Tron
,
och
den
Rättfärdighet
som
av
Tron
kommer
,
är
dess
förinnan
undertryckt
bliven
.

Men
nu
var
icke
det
yrkat
och
drivet
,
att
Bispen
deras
Herredöme
skall
bli
ifrån
tagit
,
utan
detta
allena
blir
begärt
,
att
de
vill
lida
Evangelium
må
bli
rent
predikat
och
förkunnat
,
och
att
de
vill
lösgiva
några
få
stadgar
,
vilka
utan
synd
icke
hållas
kunna
.

Likväl
till
att
undvika
vidlyftighet
,
har
vi
allena
,
de
förnämligaste
författat
,
av
vilka
man
om
de
andra
,
lättliga
kan
döma
.

Borgmästare
och
Rådmän
för
sig
och
hela
Menigheten
.

Anno
Domini
1527
.
om
Helga
Trefaldighets
tid
vi
med
vårt
älskliga
menige
Sveriges
Rikes
Råd
/
Friborne
/
Frälsemän
utan
Råds
/
Köpstadsmän
/
Bergsmän
/
och
några
fullmyndiga
bönder
utav
varje
lagsaga
kring
om
att
Riket
på
allas
deras
vägnar
som
hemma
vore
/
blir
all
denne
epters:ne
framsättningar
/
ärende
/
svar
och
beslut
/
belevade
med
alla
deras
samtycke
.

Sedan
när
då
Gud
gav
nåden
där
till
/
att
h
.
N
.
fick
så
mycket
ondarum
för
fienderna
och
tillfälle
/
var
tillhopa
kalla
Riksens
Råd
och
Adeln
som
på
den
tid
(
Gud
bättre
)
ganska
ringa
var
/
kallade
h
.
N
.
dem
tillhopa
i
Watzstena
/
och
där
bjöd
han
dem
Hövitsmans
dömt
upp
igen
/
om
de
hade
funnit
någon
god
man
där
till
fallen
hade
varit
/
och
det
hade
velat
anamma
/
och
var
överbödig
vara
honom
hörig
och
lydig
och
vaga
liv
och
hals
med
honom
för
Riket
/
ju
så
ytterligare
där
efter
som
han
rade
tillförne
begynt
hade
.

Då
nu
så
när
kom
att
landet
var
i
det
nästa
betäckt
igen
och
Stockholms
stad
skulle
uppgivas
/
fulle
I
alla
både
Ridderskapet
och
den
mene
man
till
h
.
N
.
i
Strengnes
och
bad
att
han
skulle
bli
hårda
vid
regementet
och
stå
än
nu
i
manstad
som
tillförne
Ni
ville
göra
h
.
N
.
allt
bistånd
med
liv
och
makt
/
där
skulle
han
låta
sig
uppå
så
nu
som
tillförne
/
och
till
yttermera
skäl
sade
Ni
vilja
honom
ha
för
Herre
och
Konung
över
allt
Sveriges
Rike
och
gick
strax
till
h
.
N
utväljelse
efter
Lagboken
som
han
och
då
i
de
helga
Trefaldighets
namn
där
utvalt
vart
.

Sakerna
därtill
har
h
.
N
.
väl
många
.

Och
tackar
h
.
N
.
de
Danemän
alla
mest
kring
om
att
Riket
som
här
utinnan
har
låtit
sig
finna
välvilliga
/
att
h
.
N
.
och
Riksens
Råd
icke
skulle
bli
ordlösa
män
i
Tyska
städer
/
vilka
de
har
givit
sitt
brev
och
Insegel
på
samma
gälds
betalning
/
ändå
Dalerna
allenast
dess
intet
lägga
på
hjärtat
/
utan
mena
med
uppresning
vilja
truffa
sig
till
frihet
mera
än
andra
goda
män
i
Riket
/
och
göra
andra
omlaga
med
sig
och
ha
tesliges
somliga
av
dem
givit
denna
deras
mening
så
ut
/
att
var
de
singe
den
frihet
skulle
de
väl
stillas
/
vilket
h
.
N
.
betröstar
sig
icke
till
att
inröma
dem
utan
Riksens
Råds
Råd
och
menemans
samtycke
/
som
redo
utlagt
hade
/
att
man
skulle
icke
mer
göra
dem
efter
och
egna
än
dem
i
Dalarna
/
och
sätter
det
än
nu
in
för
Er
gode
män
alla
menige
Sveriges
inbyggare
/
att
ni
ville
säga
vad
Er
där
om
synes
.

Är
och
nu
här
de
Tyska
Sändebud
till
städes
som
efter
för:ne
gälds
betalning
utsända
är
/
må
de
gode
män
av
Dalarna
och
andra
som
sig
vilja
undandraga
nu
själva
handla
med
dem
/
och
se
till
om
de
vilja
vara
betalade
med
uppresning
eller
ej
.

Sammalunda
ropas
och
emot
h
.
N
.
om
de
Borgarläge
som
han
lagt
har
i
städerna
/
Kloster
.
etc.
är
tillförne
förtäljt
att
efter
den
läglighet
på
färde
varit
har
med
detta
K
.
etc.
ärlig
/
det
vi
icke
en
alldeles
kvitte
är
/
har
nöden
tillsagt
/
att
man
skall
hålla
mera
folk
än
vant
är
/
och
tesliges
hester
/
att
de
redo
är
när
behov
görs
:
var
Gud
ville
giva
Rikena
större
säkerhet
och
rolighet
/
ville
h
.
N
.
nödigt
någon
förtunga
antingen
med
borgarläge
eller
annan
del
/
där
förinnan
säger
nöden
till
att
man
de
borgarläge
håller
/
Riksens
ränta
vill
eljest
icke
räcka
till
att
uppehålla
/
som
framledes
väl
skall
vara
förtäljt
.

Har
och
h
.
N
.
samma
predikare
en
part
här
tillstädes
och
vilja
vara
till
svars
om
deras
lärdom
om
han
är
rätt
eller
orätt
/
och
begär
att
det
måtte
ske
i
allas
Ers
närvaro
att
den
parten
som
rätt
har
må
vid
makt
bli
och
styrkas
av
alla
och
där
med
all
slik
tvedräkt
avläggas
.

Sammalunda
är
och
Kronan
försvagat
där
med
att
var
vill
vara
Konung
över
sina
egna
landbor
/
tullen
är
borta
/
Kopparberget
och
Silverberget
intet
vid
makt
/
vilket
intet
litet
avslag
är
i
Kronans
räntor
.

Kan
och
h
.
N
.
väl
besinna
att
främmande
Herrar
som
till
Riket
åstunda
/
när
de
höra
att
Svenska
män
har
sådant
sinne
att
de
är
så
lätta
på
tygeln
och
låter
sig
snarliga
förstöra
/
kunna
de
väl
snarliga
med
en
föga
kostnad
låta
här
inkomma
sådant
rykte
/
rop
och
anskre
som
de
är
redebogne
efter
löpe
att
när
i
sådan
måtte
tvedräkten
uppkommen
är
här
inbördes
/
må
de
bjuda
sig
här
till
Riket
/
som
ofta
tillförne
skett
är
:
väl
vetandes
att
all
den
stund
Sveriges
Rike
är
endräktigt
är
dem
icke
väl
möjligt
sådant
tillbedja
/
och
därför
är
det
Svenska
mannen
egen
skuld
att
här
så
ofta
har
främmande
Herrar
inkommit
och
fördärvat
Riket
/
och
därför
kan
ingen
Riksens
Herre
veta
sig
någon
trygghet
/
varken
för
utländska
eller
inländska
.

h
.
N
.
tager
den
saköre
och
fordring
som
Biskoparna
pläga
taga
att
fattiga
allmogen
icke
skall
vara
under
tu
Herrskap
.

Om
Kronans
räntor
och
Riddarskapet
som
försvagat
är
.
etc.
veta
Köpstadsmän
och
Bergsmän
ej
annat
råd
/
utan
såsom
Kyrkor
och
Kloster
har
försvagat
dem
/
så
måste
och
de
upprätta
dem
igen
/
men
hur
det
tillgå
skall
/
sätta
de
in
till
h
.
N
.
och
h
.
N:des
ärlige
Riksens
Råd
som
ena
lämpa
där
utinnan
bäst
besinna
kunna
.

Skulle
inga
Biskopar
ha
sitt
bud
till
Rohm
efter
deras
konfirmation
efter
denne
dag
.

Dessa
är
den
menemans
Svar
på
några
framsättningar
/
som
vår
nådigaste
Herre
dem
föregivit
har
,
etc.
Först
om
denne
uppstötningar
/
uppror
och
obestånd
som
årliga
års
mer
och
mer
stämplas
och
uppspringer
här
i
Riket
emot
vår
nådigaste
Herre
/
känner
Gud
att
det
är
oss
fattiga
män
ganska
lätt
att
något
sådant
företagas
skall
här
in
uti
Riket
/
emot
det
hulskap
/
troskap
och
manskap
som
h
.
N
.
lovat
vart
/
den
tid
h
.
N
.
blev
först
anammad
/
utvalt
och
utkorat
för
vår
och
Riksens
Herre
och
Konung
/
ej
allenast
då
/
utan
jämväl
i
alla
samkväm
och
Herramöte
/
vilket
den
menige
man
med
varken
med
råd
/
vet
eller
tillstärkning
oskatt
kommit
har
/
ändock
att
några
förrädare
emot
deras
ed
/
ära
och
rådlighet
begynner
något
obestånd
här
in
Rikes
/
har
dock
den
meneman
ingen
skuld
där
utinnan
/
utan
vill
heller
gärna
obrottliga
hålla
h
.
N
.
den
huldskap
/
troskap
/
manskap
som
vi
honom
lovat
och
tillsagt
har
/
viljandes
vara
h
.
N
.
hörige
/
lydige
/
hulle
och
trogne
och
stå
fasta
med
h
.
N
.
med
liv
och
makt
/
både
i
en
måtte
och
andra
/
var
behov
görs
/
och
begär
för
den
skuld
att
h
.
N
.
ville
hålla
oss
vid
lag
och
rätta
och
goda
gamla
sedvänjor
/
ville
vi
och
allesammans
vari
sin
stad
vara
allvarliga
förtänkte
att
näpsa
och
straffa
dem
som
efter
denna
dag
var
beslagen
med
förräderi
eller
obestånd
/
antingen
med
tal
eller
gärningar
emot
h
.
N
.
vare
sig
vem
det
kan
/
lekt
eller
lärt
/
tesliges
ville
vi
gärna
tillhjälpa
efter
vår
yttersta
makt
att
de
förrädare
(
som
detta
uppror
det
nu
för
hand
är
ostad
kommit
ha
)
måtte
bli
rätteligen
straffade
/
och
vem
de
helst
vara
kunna
/
och
vilja
alla
gärna
på
meniga
Sveriges
Rikes
vägnar
nu
samfälleliga
med
h
.
N
.
giva
oss
tid
upp
i
Dalarna
/
och
med
liv
och
makt
tillhjälpa
att
straffa
de
förrädare
som
detta
obestånd
ha
styrkt
och
fullföljt
/
var
h
.
N
.
oss
anders
behov
har
.

Där
näst
efter
det
att
många
munkar
(
som
fara
städse
kring
om
Riket
och
tigga
)
pläga
före
många
fåfäng
och
lögnaktig
kände
ibland
allmogen
av
vilket
den
meneman
bedragen
blir
/
enander
så
i
sanning
vara
som
de
dem
föregiva
/
genom
vilket
och
annat
sådant
förmodandes
är
/
att
sådana
uppror
eller
uppstötningar
har
endeles
sitt
ursprung
.

Tycker
oss
för
den
skuld
likt
vara
/
att
de
blir
hemma
i
deras
Kloster
/
vaktandes
de
tingest
som
dem
bör
till
Guds
tjänsten
/
dock
att
de
eller
deras
prokurator
må
utfara
två
resor
om
året
/
en
om
sommaren
annan
om
vintern
/
efter
deras
näring
var
resa
icke
längre
ute
än
en
månad
.

Yttermera
som
h
.
N
.
berör
om
de
borglige
/
har
den
meneman
alldeles
intet
där
om
talat
/
varken
lönnligen
eller
uppenbarligen
efter
det
rör
oss
intet
an
/
utan
tycker
oss
väl
likt
vara
/
att
Klostren
hålla
borgarläge
/
vart
efter
som
det
har
makt
till
/
dock
är
tillbörligt
/
att
där
måtte
skickas
gode
karlar
till
Klostren
/
som
utan
all
buller
eller
skalkhet
sig
med
späkt
har
kunnat
låtandes
sig
åtnöja
med
den
del
som
de
fattiga
män
har
att
skifta
med
dem
/
och
att
de
icke
heller
gör
något
övervåld
som
där
omkring
Klostren
bo
/
sammaledes
att
Guds
lidgård
icke
förhindras
i
Klostren
någraledes
.

Om
de
andra
artiklar
där
vi
icke
kunde
svara
till
/
som
är
om
Kyrkans
räntor
och
andra
sådana
sätter
vi
in
till
vår
K
.
N
.
Herre
och
Riksens
Råd
.
etc.
ganska
högliga
och
ödmjuka
bedjandes
Ers
Nåds
Högmäktighet
.

Vi
efterskrivna
Johan
med
Guds
nåd
Greve
till
Hoghn
Brockenhusen
.
etc.
Hövitsman
på
Wijborgh
.
etc.
Ture
Jönson
Riddare
vår
nådigaste
Herres
Hovmästare
/
Lars
Siggeßon
Marsk
/
Holger
Carson
Riddare
/
Axell
Påße
/
Michell
Nilßon
Laghman
/
Nils
Olßon
/
Iffuar
Flämingh
/
Axell
Anderßon
/
Knut
Anderßon
/
Nils
Claußon
/
Jord
Bonde
/
Pedher
Hanßon
/
Biorn
Claußon
/
Hendrich
Ärlanßon
/
Pädher
Ärlaßon
Sveriges
Rikes
Råd
.
etc.
Gör
vitterligt
/
att
som
vi
här
församlade
var
i
Westerårs
efter
vår
nådige
Herres
Konung
Göstaffz
skrivelse
med
menige
frälset
av
allt
landet
/
tesliges
Köpstadsmän
/
bergsmän
och
några
fullmunniga
av
varje
Lagsaga
kring
om
allt
Riket
:

Gav
samme
vår
nådige
Herre
oss
förre
några
märkliga
brister
som
i
Riket
vore
/
varför
han
ingalunda
betrösta
sig
längrr
bli
vid
Riksens
regemente
och
styrelse
med
mindre
samma
brister
botade
var
:
och
bad
oss
alla
samman
brister
överväga
och
finna
där
råd
emot
/
annars
ville
han
uppsäga
oss
Riket
igen
/
att
vi
där
om
besörjde
det
bästa
vi
kunde
/
ibland
vilka
brister
våra
denna
de
yppersta
de
och
väl
så
viktiga
vore
/
att
de
väl
måtte
göra
en
vederstyggelse
vid
Riksens
Regemente
/
som
Hans
Nåd
och
somliga
av
dem
hade
allaredan
tillförne
föregivit
/
då
han
vart
utkorad
för
Herre
och
Konung
över
Riket
.

Den
tredje
bristen
var
att
h
.
Nåds
Riddarskap
var
svarliga
försvagad
och
behövde
för
den
skull
alltid
bedjas
hjälp
av
Kronan
(
som
intet
under
vår
)
och
var
Kronans
del
desto
mindre
för
Konungens
uppehälle
.

Fjärde
brist
/
att
Hans
Nåd
påfördes
mångestädes
i
Riket
att
han
låter
indraga
nya
tro
/
och
att
det
mest
gjorde
en
stor
del
av
präster
och
munkar
/
därför
att
h
.
Nåd
kunde
lida
dem
som
predikade
rena
Guds
ord
och
Evangelium
det
de
icke
höra
eller
lida
måtte
.

Till
att
bota
den
andra
/
säger
vi
att
efter
den
ränta
/
som
Bisperna
/
Domkyrkorna
/
Kaniker
/
och
Kloster
har
/
är
kommen
från
Riksens
inbyggare
och
med
Herrarnas
stadfästelse
som
då
var
;
Därför
samtycker
vi
alla
med
för:ne
vår
nådiga
Herre
/
att
Kronans
ränta
den
nu
förminskat
är
/
må
där
med
upprättas
igen
.

Därför
på
det
att
Riket
skall
vara
den
fara
för
utan
efter
denna
dag
/
samtycker
vi
alla
för
oss
/
för
våra
efterkommande
/
att
de
efter
denna
dag
icke
skulle
rida
med
/
flera
karlar
än
som
för:ne
vår
nådiga
Herre
dem
föresäger
.

Vad
över
är
i
deras
uppbörd
det
kommer
till
att
föröka
Kronans
ränta
där
med
så
att
de
skulle
giva
Konungen
ett
stycke
penningar
/
efter
som
de
kunna
med
honom
över
ens
vara
/
och
där
till
antvarda
honom
de
Slott
och
fästen
som
de
nu
har
.

Sammalunda
ske
med
Domkyrkornas
och
Kanikernas
ränta
/
när
överlagt
är
vad
till
deras
redliga
uppehälle
behövs
/
då
tar
Konungen
det
utöver
är
/
i
deras
ränta
/
uti
ett
stycke
penningar
sig
till
hjälpa
.

Samtycker
vi
att
här
efter
skicka
Konungen
en
god
Riddarmans
man
utöver
samma
Kloster
den
Klosterfolket
skall
låta
få
sitt
redliga
uppehälle
och
Klostret
vid
makt
håller
/
vad
där
utöver
kan
vara
/
gör
han
Konungen
tjänst
utav
med
borgarlägga
eller
eljest
som
Konungen
täckes
.

Och
som
Gud
förbjuda
att
någon
skada
eller
fördärv
hända
för
för:na
handel
skull
i
Riket
på
vår
Nådiga
Herre
eller
någon
av
oss
utav
inländska
eller
utländska
;
Bepliktar
vi
oss
först
med
vår
nådiga
Herre
/
att
var
och
en
utav
oss
samma
skada
och
fördärv
avvärja
med
liv
och
makt
;
yttermera
om
någon
utav
oss
antingen
innan
rads
eller
utan
/
ädla
eller
oädla
/
Köpstadsman
eller
bonde
sig
härifrån
sins
drar
och
förmärkt
blir
med
tal
/
ord
eller
gärningar
/
lönnliga
eller
uppenbarliga
/
den
ville
vi
för:de
Sveriges
Rikes
Råd
/
frälsemän
/
Köpstadsmän
/
Borgmästare
och
den
menige
mans
fullmyndige
av
varje
lagsaga
/
tillhjälpa
att
han
straffas
skall
.

Och
har
vi
här
med
vårt
Riksens
Råd
och
tesliges
med
menige
frälset
/
Köpstadsmän
/
Bergsmän
och
mene
Allmogens
fullmyndiga
Sändebud
näst
Guds
hjälp
övervägt
allas
Ers
bästa
och
långliga
bestånd
/
som
Ni
väl
förnimmandes
var
/
uti
Riksens
Råds
brev
/
som
här
med
följer
och
förste
vi
oss
fulleliga
till
Er
alla
/
att
vi
Er
alltid
ha
skulle
för
tro
och
välvilliga
undersåtar
/
vi
ville
däremot
för
Er
och
alla
Sveriges
Inbyggares
bästa
/
ha
ospard
var
hals
och
välfärd
/
där
må
i
Er
alla
fulleliga
på
förlåta
/
vad
yttermera
förhandlat
och
beslutat
blev
i
för:ne
möte
/
kunde
denne
er
fullmyndiga
Sändebud
själva
giva
er
tillkänna
.

Riksens
Råds
Brev
till
den
meneman
.

Biskopar
vi
ingen
till
Präster
/
utan
den
som
kan
predika
för
Folket
Guds
Ord
.

Prelaturer
/
Canonier
och
Prebender
/
skola
ej
förses
med
mindre
Konungen
blir
åtspord
/
eller
den
hans
Nåd
där
till
skickandes
var
.

Händer
Fästman
lägra
sina
Piga
eller
Lagfästa
Hustru
/
bötar
där
intet
före
/
efter
emellan
dem
är
rätt
Äktenskap
för
Gud
/
och
må
han
icke
åtskiljas
vid
henne
.

Överger
han
henne
/
straffas
efter
Lagen
.

Icke
skall
heller
något
sjukt
Folk
tvingas
av
Prästerna
till
något
Testamente
emot
deras
fria
Vilja
.

Ingen
uppehåller
Sakramentet
för
några
om
Påsk
eller
annan
Tid
/
antingen
för
Gäld
eller
annat
/
utan
söker
Präster
och
Kyrkor
sin
rätt
på
Ting
och
Stämma
/
som
förberört
är
.

Svarade
Nils
att
han
hade
(
misstankar
till
)
honom
,
att
han
skall
ha
burit
det
bort
i
Ölsmål
,
(
efter
han
en
gång
tillförne
hade
burit
bort
ett
stop
i
Ölsmål
,
)
(
Så
medan
det
var
allenast
en
misstanke
vart
sagt
att
de
skulle
förlikas
medan
det
var
i
hastiga
mod
skett
,
då
sade
Morthen
att
han
ville
göra
sig
därför
själv
tolfte
fri
och
Lade
fram
deras
handskar
som
hade
lovat
gå
med
sig
,
Så
medan
det
var
en
misstanke
och
skedde
med
hastigt
mod
vart
förlikat
och
lades
40
daler
i
vite
den
Morthen
därför
förviter
.
)
Morthen
kärade
till
Nils
Höös
om
(
en
del
i
)
en
Brännvins
Panna
,
vart
sagt
att
Nils
skulle
giva
där
för
2
mr
Penningar
.

Den
12
December
höll
högbetrodd
Jahan
Jacobsson
Kamrer
(
och
Häradshövding
)
Lagting
uti
Befallningsmannens
Ädel
och
välbördig
Albrecht
Magduwals
närvaro
dessa
Edsvurna
såtar
i
Nämnden
.

Då
svarade
Allmogen
,
att
Fogden
och
Skrivaren
har
nog
där
på
drivit
,
men
för
det
att
föret
slog
så
hastigt
av
och
en
del
för
stor
fattigdom
icke
komma
fram
,
det
är
orsaken
,
då
förmanades
dem
som
är
tillbaka
att
de
Låta
komma
fram
till
bruket
det
de
skyldiga
är
vid
bot
.
)
h
.
Elin
i
Bokarby
lät
förste
sin
uppbjuda
sitt
hemman
som
Olof
Andersson
hade
tagit
av
henne
till
köps
och
givit
henne
därpå
12
lod
silver
lodet
för
2
mr
och
10
daler
Penningar
då
tillfrågades
Olof
Nilsson
hennes
Son
om
han
icke
ville
behålla
.

Så
hade
han
och
givit
alla
dessa
förarna
tillhopa
i
vängåvor
eller
Stille
Penningar
4
daler
.

Item
hade
fönne
Staphan
köpt
av
h
.
Christin
Per
Nilssons
i
Akra
ett
öres
Land
Jord
och
husen
och
givit
henne
därför
472
daler
Penningar
.

Item
hade
han
slagit
Morthens
Piga
en
Pust
vart
därför
sak
3
mr
.

Olof
i
Bengzbo
,
Giesmyre
och
Fänebeckiekarlarna
kärade
att
Matz
i
Långrudhe
hade
stänkt
allt
för
mycket
skog
in
.

Staphan
i
Hof
är
kommen
i
rykte
för
sin
lege
Piga
,
och
är
han
skylld
samma
jänta
då
bekände
Staphan
att
han
Låg
när
henne
en
natt
,
men
fönne
Brita
som
är
belägrat
av
Staphans
dräng
Hans
,
sade
att
hon
Låg
hos
honom
tre
nätter
åt
slag
i
en
vecka
,
Staphan
fäste
Lag
att
göra
sig
fri
själv
12
nästa
ting
.

Vart
för
den
skull
han
sak
80
daler
och
hon
40
daler
på
h
.
M:ttz
Drottningens
nådiga
behag
.

Vart
förenade
och
Lades
20
daler
i
vi
de
den
sig
på
den
andra
först
förbryter
.

Anders
Skomakare
hade
gått
objuden
till
gästbod
vart
sak
3
mr
.

Vart
sak
3
mr
för
vardera
Hans
i
Libbarebo
hade
brutit
det
vi
de
som
är
satt
emellan
honom
och
hans
granne
år
1619
den
10
Martij
(
N.3
)
40
mr
.

Bekom
och
Pers
hustru
Syster
Penningar
av
Erich
Olofsson
,
och
fördenskull
har
M
.
Jöran
intet
henne
tilltala
)
Anders
Perssons
hustru
Syster
i
Göthebrunna
Elin
Anders
dotter
stod
in
för
rätten
och
till
stod
sig
ha
uppburit
av
h
.
Karin
Erich
Abramssons
i
Hökeby
medan
hon
var
Änka
Penning
10
daler
(
,
vilka
Penningar
hon
bekom
i
Skärplinge
i
Löfsta
Socken
av
Erich
Brom
för
sitt
möderne
och
Lade
dem
ned
i
Hökeby
.
varför
Elin
Andersdotter
avhände
sig
och
sina
efterkommande
och
till
ägnade
2
)
h
.
Karin
och
hennes
arvingar
till
evärdlig
egendom
.

Matz
Benchtsson
i
Långerudhe
och
Thomas
Matsson
i
Läby
i
Börklinge
Socken
och
deras
bröder
och
Systrar
har
uppburit
av
S
.
Olof
skrivare
Penningar
7
daler
.
(
Item
har
de
uppburit
att
h
.
Karin
Penningar
17
daler
.

Michil
Olofsson
i
Karby
berättade
att
Jöran
Crutz
borgare
i
Gäfle
hade
sänt
till
honom
25
få
Torra
gäddor
och
Abborrar
Smör
18
mr
och
en
halv
tunna
Lax
näst
för
Julen
hade
fönne
Michil
begärt
lov
av
HäradsFogden
att
sälja
samma
fisk
det
han
och
lovade
,
dock
sedan
han
förnam
att
han
hade
*
sålt
något
där
av
till
8
få
.
av
vilka
8
få
Erich
Olofsson
tog
5
få
efter
sitt
Betzman
och
ändå
kastat
bort
vidjorna
som
de
vore
ombundna
med
,
då
tog
Erich
Olofsson
ifrån
honom
17
få
Tonfisk
.

Thomas
i
Grytteby
Per
Larsson
i
Bolmyra
lät
tredje
sin
uppbjuda
2
öres
Land
Jord
och
hus
som
han
köpt
hade
av
Morthen
Larsson
Ryttare
och
hans
Systrar
Barbara
och
Malin
Lars
döttrar
(
för
16
daler
Pegr
och
en
spann
vete
i
Stille
Item
gav
han
Thomas
i
Grytheby
i
Stille
eller
vänskapsgåvor
en
treggie
lod
silver
sked
efter
han
är
i
börden
)
.

Anders
Persson
i
Göthebrunna
stod
här
och
lov
gav
(
h
.
Karin
S
.
Erich
Abramssons
på
sin
barns
vägnar
att
lossa
av
honom
sin
del
i
Hökeby
)
där
på
han
räckte
Anders
Höök
handen
efter
han
är
barnens
Målsman
.

Ma:ttz
Befallningsmans
Ärlig
och
välbetrodd
Hans
Jönssons
närvaro
,
dessa
Edsvurna
såtar
i
Nämnden
.

Item
hade
hennes
barns
fäder
fader
Hans
Andersson
köpt
av
Erich
Larsson
i
Vpsala
någon
Jord
som
köpebrevet
vidare
utvisar
.

Vad
Katzlinge
vidkommer
som
Michil
Morthess
hade
bort
bytt
för
Myrkarsbo
för
24
år
sedan
hade
varken
i
hans
livstid
eller
sedan
han
död
blev
,
varit
Klandrat
för
än
nu
detta
år
624
av
hans
måg
som
på
Myrkarsbo
bor
såsom
och
hans
Son
som
än
i
livet
är
,
vilka
för
menar
sig
vilja
göra
bytet
om
intet
som
emellan
deras
fader
Michil
Morthensson
och
Anders
Erichsson
,
efter
där
med
icke
är
Lagligen
tillgånget
som
uti
det
10
Kap.
i
Jorda
Balken
står
förmält
.

Lasse
Andersson
i
Westerekeby
hade
dolt
en
liten
kille
som
var
kommen
in
i
hans
gård
och
intet
upplyst
den
vart
sak
3
mr
Lades
vite
40
mr
att
ingen
må
förvita
honom
därför
.

Olof
Persson
i
Laghmyra
hade
tagit
en
Yxa
olovandes
på
vägen
av
Michil
Erchsson
i
Granby
i
Börklinge
vart
sak
6
mr
.

Pedher
Anderson
i
Smedby
var
Stämd
att
Svara
Arrendatorn
,
vart
Saker
till
3
.
mr
.
till
vidare
Rannsakning
.

Men
där
han
här
efter
övergiver
henne
skulle
han
vara
saker
till
40
.
mr
.

Och
sedan
be:te
Lars
Jönsson
var
Förrymd
hade
Erich
Pedersson
bortdolt
Älghuden
och
henne
gömt
Under
sitt
Stuggolv
,
där
Läns
och
Fjärdings
Mannen
sedan
hade
Funnit
henne
Igen
,
och
Allden
Stund
be:te
Erich
Pedersson
hade
Uti
Sanning
dolt
och
gömt
med
be:te
Larss
Jönsson
,
därför
var
han
Lika
delaktig
med
be:te
Larss
Jönsson
Uti
Saken
kunde
För
den
skull
Nämnden
Icke
Fria
honom
Ifrån
den
dom
Som
Hans
Konung
Ma:tz
Brev
Innehåller
,
Blev
därför
be:te
Erich
Pederssonn
sagt
att
föras
över
med
bo
och
bohag
till
Jngermanne
Land
.

Sedan
Hade
be:te
Erich
OluffSon
Slagit
be:te
Pelle
Pederssonn
igen
tre
blånader
med
en
Stor
,
där
till
han
ej
Nekade
Utan
sade
att
han
måtte
något
tagas
till
och
värja
sig
med
,
vart
därför
Saker
till
9
mr
.

Hans
Jörnssonn
i
väster
Ekeby
var
stämd
av
Nämnde
Mannen
,
att
Svara
Arrendatorn
vart
saker
till
3
mr
för
Svarlösa
till
vidare
,
rannsakning
.

Morthen
i
Torkilsbo
hade
klagomål
på
sig
var
stämd
kom
intet
vart
sak
3
mr
.

Kärade
och
Anders
Andersson
Höök
Länsman
att
hans
S
.
fader
Anders
Hock
Häradsskrivare
hade
betalat
Kronan
en
stor
hop
för
Holfwebo
hemmanet
som
(
han
framledes
bevisa
ville
)
.

Noch
Hans
broder
som
kniven
drog
till
att
göra
skada
,
dock
ingen
gjorde
,
Sakfälldes
till
Penningar
—
3
mr
.

Noch
vittnade
Nämndemännen
samt
andra
inhäradsmän
,
att
Ädle
och
välbördig
Magduualtz
bönder
,
är
så
väl
de
,
såsom
hans
Sättegårdh
Uti
en
Boollby
,
N
:

Till
vilket
be:te
Duwalt
och
sade
sig
Lika
Såsom
han
Arrendet
av
Hennes
M:tz
S
.
och
höglovlig
åminnelse
först
fångat
har
,
med
Utsäde
av
gamla
Rågen
Levererat
.

Nottegarn
,
vilka
han
av
Tijerph
Socken
på
Petters
år
Uppburit
hade
,
det
Hans
Jönsson
icke
heller
Neka
kunde
:

Noch
vittnade
Nämndemännen
samt
andra
inhärads
män
att
Hoffqwarn
,
har
av
ålder
Lytt
och
Legat
Under
Örby
gård
,
är
och
Upprättat
med
Örby
Läns
omkostnad
.

Be:te
Horkona
brijta
anders
dotter
är
tillförne
dömd
,
och
Utav
den
höglovlige
Kung:
Hovrätten
till
bötet
40
dr
resolverat
.

Och
vad
mera
hennes
S
.
svärfaders
gäld
ännu
Restera
kunde
,
avdömdes
att
alla
Arvingarna
skola
där
om
Lika
delaktiga
vara
,
var
och
en
efter
den
kvota
de
ärvt
har
.

Därnäst
företogs
följande
uppbud
och
intäckningar
.

Ävenledes
blev
på
Gustaf
Michelssons
anhållan
skatte
och
besittnings
rätten
av
bemälda
hemman
i
ÖsterEkeby
honom
,
Gustaf
Michelsson
,
till
handa
tredje
gången
uppbjuden
till
följe
av
bytes
brevet
,
som
så
väl
nu
som
vid
förra
tinget
uppvisat
och
uppläst
blev
.

Kronobefallningsmannen
välbetrodde
Petter
Yckenberg
lät
uppläsa
högvälborne
herr
baron
och
landshövdingens
brev
och
ordres
till
sig
av
den
23
maj
sistlidne
angående
förenings
träffande
om
en
viss
brandstods
utgörande
hädan
efter
,
likmätigt
Kungl.
Maij:t
därom
till
högvälbemälda
herre
avlåtna
nådigaste
/
brev
och
skrivelse
av
den
28
martij
sistlidne
,
begärandes
herr
befallningsmannen
,
det
ville
socknens
förmodligen
utsedde
fullmäktige
yttra
sin
mening
därom
.

Eljest
hade
han
också
instämt
Michel
Andersson
,
för
det
han
hela
nästlidet
år
försummat
att
prestera
sin
hållskjuts
vid
gästgivare
gården
,
vilken
emedan
han
där
till
intet
neka
kunde
utan
sade
,
att
Swen
Pärsson
i
Tårkelsbo
är
orsaken
där
till
,
som
lovat
skjutsa
för
honom
men
det
intet
hållit
;
Ty
prövas
skäligt
,
det
bör
Michel
Andersson
för
en
slik
hållskjuts
eftersättande
böta
sina
3
gånger
3
marker
silvermynt
efter
1664
års
gästgivareordnings
13
§
,
kunnandes
han
söka
Swen
Pärsson
igen
,
om
han
gitter
och
förmenar
sig
ha
skäl
där
till
.

Annicka
Erichsdotter
nekade
härtill
och
sade
,
att
hon
intet
sänglag
haft
med
Petter
Silfverdahl
.

åter
igen
Erich
Pärsson
i
Labärga
angående
den
väg
,
varom
de
vid
sista
ting
tvistade
,
med
påstående
,
det
måtte
han
antingen
få
bemälda
väg
fram
emellan
Huusby
fjäll
i
Karby
gärde
och
Labärga
äng
,
såsom
han
i
förra
tider
gått
,
och
att
Erich
Pärsson
till
den
ändan
skall
böra
taga
upp
sin
gärdesgård
och
flytta
honom
längre
in
åt
,
/
därest
han
till
förene
stått
,
eller
och
låta
honom
,
efter
senare
tiders
överenskommelse
,
ha
vägen
över
Labärga
äng
i
stället
.
2:do
expenser
efter
räkning
till
13
daler
30
.
/
.
kopparmynt
.

Erich
Pärsson
sade
sig
intet
kunna
svara
här
till
,
efter
som
hemmanet
intet
hör
honom
utan
dess
stugbarn
till
,
varför
han
menade
,
det
deras
målsmän
eller
förmyndare
böra
härom
stämmas
och
höras
,
innan
något
visst
härom
slutas
kan
.

Men
på
rättens
/
interposition
gav
Erich
Pärsson
äntligen
Olof
Olssön
den
oförrätt
han
gjort
honom
medelst
berörda
skimpfelige
expressioner
,
som
förra
protokollet
vid
handen
ger
,
efter
som
Olof
Olssön
bad
honom
om
förlåtelse
och
tillstod
,
att
det
skedde
av
ett
hastigt
överilande
,
men
expenser
ville
Erich
lika
fullt
ha
av
Olof
.

Mårten
Mattsson
i
Allerbäcke
och
Johan
Olssön
i
Grytby
hade
var
annan
instämt
,
den
förra
den
senare
angående
det
Johan
Olssön
skall
uppå
en
av
honom
presenterad
obligation
begärt
och
fått
uppbjöd
å
Mårten
Mattssons
hemman
i
Allerbäcke
,
det
han
så
mycket
mera
vill
ogilla
och
har
upphävit
,
som
han
aldrig
skall
utgivit
en
slik
obligation
eller
sätt
sitt
namn
och
bomärke
därunder
,
mycket
mindre
det
bomärke
,
som
/
står
under
obligationen
,
emedan
han
aldrig
skall
brukat
ett
sådant
bomärke
,
viljandes
fördenskull
,
det
Johan
Olssön
skall
bevisa
,
att
han
givit
en
slik
obligation
ifrån
sig
och
sätt
bomärket
därunder
,
eller
bli
därför
efter
lag
ansedd
,
så
väl
som
för
det
han
skall
betingat
sig
för
stort
intresse
,
nämligen
i
tunna
.
säd
om
året
för
lånet
av
180
daler
'
kopparmynt
;
den
senare
den
förra
med
påstående
,
att
Mårten
Mattsson
själv
kommit
till
honom
med
obligationen
och
själv
ritat
bomärket
därunder
uti
Johan
Olssons
stuga
,
vilket
ock
så
mycket
mera
skall
kunna
finnas
och
slutas
vara
sant
,
som
han
intet
skall
kunnat
,
utan
revers
och
behörig
säkerhet
av
hemmanets
pantsätttande
,
låna
honom
,
såsom
då
för
tiden
,
nämligen
år
1720
,
när
lånet
gjordes
till
hemmanets
skatterättighets
lösen
ifrån
Kungl.
Maij:tt
och
Kronan
,
varande
en
lös
och
ledig
dräng
,
beklagandes
,
att
han
med
en
sådan
otack
och
skamlig
tillvitelse
skall
bli
bemött
för
sin
honom
gjorde
välgärning
,
helst
han
intet
betingat
sig
ovanberövade
intresse
utan
tagit
obligationen
sådan
emot
,
som
han
var
skriven
,
till
bevis
att
han
borde
ha
för
/
skrivit
intresse
av
Mårten
Mattsson
för
sitt
gjorda
lån
,
viljandes
fördenskull
,
det
Mårten
Mattsson
måtte
själv
lagligen
omgälla
det
han
honom
ärnat
.

Emedan
Lars
Olssön
Brundin
såsom
hallnabrukare
av
bokhållaren
Christian
Ohsengii
skattehemman
Tälsgiärde
/
njutit
hälften
av
allt
vad
hemmanet
kastat
av
sig
och
det
,
skönt
intet
kontrakt
är
emellan
jordägaren
och
hallnabrukaren
,
ändå
alltid
är
brukligt
,
att
hallnabrukaren
svarar
till
hälften
uti
knektehållet
;
alltså
kan
tingsrätten
intet
annat
finna
,
än
att
Lars
Olssön
bör
,
efter
Ohsengii
utlåtelse
,
åtminstone
bestå
1
/
3
del
av
den
nylagde
soldatens
lön
,
lega
och
städsel
i
proportion
av
det
,
som
därav
på
Tälsgiärde
hemmanet
sig
kan
belöpa
,
efter
som
han
intet
längre
blir
vid
hemmanet
än
till
nästkommande
midfasta
.

Om
de
påstådda
forpenningarna
,
som
Lars
Olssön
nekat
sig
ha
lovat
,
och
de
2:ne
öke
dagsverken
,
som
Ohsengius
skall
fått
av
Brundin
men
den
förra
där
till
nekat
,
lämnas
dem
å
båda
sidor
att
stämma
var
annan
till
nästa
ting
och
,
om
de
gitta
,
varannan
det
överbevisa
,
efter
som
ingendera
disputerat
det
begärda
uppskovet
där
med
.

Till
följe
av
högvälborne
herr
baron
och
landshövdingens
givna
resolution
uppå
framlidne
häradsskrivarens
Petter
Agrells
efterlåtna
änkas
,
dygdesamma
hustrus
Elisabeth
Wendlers
,
supplique
undersöktes
nu
om
hennes
tillstånd
,
och
som
nämnden
med
flera
närvarande
visste
att
intyga
,
det
hon
är
en
gammal
människa
in
emot
70
år
samt
sjuklig
och
krasslig
,
utan
att
ha
någon
annan
egendom
än
1
/
2
skattefrälsehemman
,
varandes
nu
i
det
tillstånd
stadd
,
att
om
hon
intet
hade
sin
måg
,
sergeanten
äreborne
och
manhaftig
Benjamin
Elgklo
,
att
lita
sig
till
,
så
förmådde
hon
intet
att
så
sköta
och
förestå
bemälda
hemman
,
att
hon
därav
kunde
ha
sin
föda
och
utkomst
,
utan
var
i
annan
händelse
råkandes
i
uselhet
och
armod
;
Ty
blev
detta
till
bevis
därom
meddelat
.
/

S
.
T
.
Gör
här
med
veterligt
,
att
år
efter
vår
Herres
och
frälsares
Jesu
Christi
nåderika
födelse
1736
den
27
\
zxM,arii
,
då
jag
rätt
laga
ting
höll
med
allmogen
och
menige
man
av
Wendels
tingslag
på
vanligt
tingsställe
uti
Karby
by
,
när
varande
Kronans
länsman
välaktat
Gabriel
Wretberg
och
tingslagets
nedanskrivna
vanliga
nämnd
,
lät
kyrkoherden
i
Dannemora
ärevyrdige
och
högvällärde
herr
Erich
Ekeroth
anhålla
om
denna
rätts
faste
och
stadfästelse
brev
å
skatte
och
besittningsrätten
av
det
frälsehemman
i
Kläringe
,
bestående
av
7
/
8
mantal
,
vilket
frälseåboen
Pär
Hansson
innehaft
och
åbott
.

Responsum
,
i
14
år
.

brev
av
den
7
juli
1692
och
5
november
1694
,
bör
efter
orden
förstås
utan
någon
annan
uttydning
;
och
som
nästbemälda
kontrakt
förmår
och
innehåller
uti
dess
6
§
,
att
Michel
Andersson
skulle
vara
ansvarig
och
fullgöra
allt
vad
efter
det
med
herr
rådman
Almgreen
slutna
kontraktet
intet
var
fullgjort
och
efterkommit
,
samt
uti
den
7
§
,
att
han
skulle
visa
,
hur
han
använt
husrötesumman
efter
1725
års
syn
,
eller
i
brist
därav
sådant
utbetala
tillika
med
den
husröta
,
som
sedermera
kunde
vid
gården
vara
existerad
;
varandes
det
en
klar
analogi
och
likhet
,
att
om
Ahlsteen
kunde
njuta
sådant
till
godo
,
sedan
han
hade
köpt
hemmanet
av
Almgreen
,
det
Anders
Andersson
även
bör
njuta
samma
förmån
efter
Ahlsteen
.

I
annan
händelse
bör
de
vad
som
dem
,
såsom
ovanförmält
finns
,
påfört
är
,
strax
betala
eller
undergå
exekution
,
varifrån
dock
Anders
Ersson
i
Uggelbo
befrias
,
till
dess
det
efter
föregången
ytterligare
stämning
närmare
blir
bevisat
,
huruvida
han
bör
njuta
sin
uppvisade
slutsedel
till
godo
eller
intet
.

Om
de
frånvarande
kan
tingsrätten
sig
intet
utlåta
,
innan
det
visas
,
att
de
blivit
vederbörligen
/
stämde
,
som
denna
gången
intet
skett
.

För
Anders
Erssons
i
Jordansbo
,
nu
i
Åkra
,
169
daler
*
,
som
erkände
blev
,
gick
befallningsmannen
Philip5
Befwert
i
caution
,
så
att
de
inom
2
år
skulle
bli
betalda
,
och
efter
som
Lidberg
lät
sig
där
med
åtnöja
,
så
förblir
det
ock
där
vid
.

Länsmannen
Gabriel
Wretberg
anklagade
också
gifte
drängen
Nils
Pärsson
,
som
skall
vistas
hos
mjölnaränkan
i
Bergby
,
och
ladugårdspigan
hustru
Eva
på
Storgården
ibidem
,
för
det
de
nästlidne
långfredag
skola
varit
druckna
samt
kivat
och
slagits
sins
emellan
,
så
att
Nils
fått
både
blånader
och
blodviten
,
påståendes
därför
den
plikt
emot
dem
,
som
lag
förmår
.

Hustru
Eva
tillstod
,
att
allt
så
tillgått
,
som
vittnet
berättat
,
men
nekade
ännu
,
att
hon
slagit
eller
tillfogat
Nils
någon
åkomma
,
utan
lär
han
,
sade
hon
,
ha
stött
sig
,
när
han
for
efter
henne
i
mörkret
och
hof
henne
ut
ur
stugan
.

Erich
Pärsson
och
Michel
Nilsson
ville
,
efter
sin
vice
versa
stämning
,
det
denna
sak
måtte
stå
oavgjord
,
till
dess
barnen
bli
myndiga
,
att
de
själva
få
försvara
sin
rätt
,
emedan
det
intet
vill
anstå
dem
att
samtycka
till
någotdera
i
mellertid
,
efter
som
det
intet
kan
avlöpa
utan
stor
olägenhet
och
skada
för
ängen
.

Mårten
Mattsson
,
som
först
i
går
blivit
stämd
,
ville
intet
svara
,
innan
han
blir
lagligen
stämd
;
vilket
tingsrätten
,
efter
processen
,
intet
ogilla
kunde
,
utan
anstår
alltså
här
med
,
vad
honom
angår
,
till
dess
han
blir
lagligen
stämd
.

Erich
Mattsson
förnams
vara
nyss
kommen
till
hemmanet
och
har
således
intet
vetat
av
sin
hålldag
,
helst
han
icke
heller
var
till
kyrkan
den
gången
,
när
det
blev
tillsagt
om
hållskjutsen
;
varför
ock
han
från
böter
denna
gången
befriad
/
var
,
men
så
bör
han
likväl
uppfylla
denna
skjuts
,
enär
han
påkallad
var
till
gästgivare
gården
.

Ersättning
för
det
Brundin
haft
Ohsengii
häst
till
Strömsberg
med
utlagssäden
ville
han
så
mycket
mindre
bestå
,
som
han
jämwäl
då
förde
Ohsengii
egen
säd
med
.

Om
dagsverken
menade
Brundin
vara
vid
sista
ting
dömt
;
men
sina
i
|
ökedagsverken
gav
han
efter
emot
den
säd
han
fått
av
det
nyupptagna
åkerstycket
,
som
Ohs
begärt
.

Och
emedan
det
intet
kunnat
finnas
,
att
Brundin
haft
någon
ond
mening
med
det
han
lämnade
den
av
ålder
och
fodernöd
död
blivna
hästen
i
ladugården
liggande
tills
nu
i
vår
eller
att
han
i
orättan
tid
flyttat
från
hemmanet
,
efter
som
midfastan
kom
mycket
sent
i
år
,
vid
den
tiden
man
eljest
plägade
både
träda
och
så
,
så
frierkänns
han
även
därutinnan
från
Ohsengii
tilltal
.

Men
för
det
Brundin
haft
Ohsengii
häst
till
Strömsberg
med
utlagssäden
bör
han
honom
betala
,
efter
som
han
i
kontraktets
9
§
sig
förbundit
till
att
föra
den
bort
,
dock
det
allenast
med
2
daler
14
.
/
.
kopparmynt
,
emedan
Ohsengius
haft
2
fjärdingar
egen
säd
däribland
,
åliggandes
ock
honom
,
Brun
/
din
,
att
själv
bestå
kyrko
och
bogårds
byggnaden
med
de
där
till
använda
gångled
,
emedan
sådant
alltid
hör
en
hallnabrukare
till
att
göra
,
efter
som
kontraktet
emellan
honom
och
jordägaren
intet
uttryckligen
frikallar
honom
därifrån
.

Quasstio
till
länsmannen
,
när
och
varest
han
befanns
drucken
?

Responsum
,
under
högmässopredikan
uti
vapen
huset
,
därest
han
skall
funnits
av
drycker
så
betagen
,
att
han
så
när
hade
raglat
omkull
och
,
när
han
gick
ut
,
lämnade
efter
sig
både
hatt
och
käpp
,
skolandes
han
,
som
länsmannen
sade
,
intet
varit
drucken
under
ottensångspredikan
,
varav
han
menade
nogsamt
kunna
finnas
,
det
han
måtte
ha
emellan
predikningarna
varit
/
inne
på
Håfgårdzberg
hos
skolmästare
Brödernas
och
tagit
för
mycket
till
livs
antingen
av
öl
eller
brännvin
.

De
avlade
alltså
ojävade
vittneseden
och
berättade
därefter
var
för
sig
,
först
Anders
Olssön
,
att
när
gudstjänsten
till
högmässan
begyntes
,
skall
han
,
efter
han
fann
sig
något
opasslig
,
satt
sig
ute
i
vapenhuset
,
varefter
Ekeroth
skall
kommit
raglandes
in
och
satt
sig
på
skalmen
av
likbåren
samt
släppt
hatten
ifrån
sig
.

Sedan
han
där
hade
suttit
en
liten
stund
,
skall
han
gått
in
till
vapenhusdörren
och
givit
sig
till
att
se
i
bok
med
en
annan
samt
vid
detsamma
raglat
in
på
lektorn
vid
Strengnäs
gymnasium
herr
magister
Stenius
,
som
då
stod
där
vid
dörren
,
så
att
han
måste
vika
undan
för
honom
,
varefter
Ekeroth
skall
gått
raglandes
tillbaka
till
båren
och
äntligen
gått
därifrån
ut
,
lämnandes
både
hatt
och
käpp
efter
sig
,
varför
han
med
flera
,
som
stod
i
vapenhuset
den
gången
,
skola
bett
Olof
Larsson
taga
upp
hans
hatt
och
käpp
och
gå
ut
till
honom
med
samt
bedja
honom
,
till
vidare
förargelses
förekommande
,
bli
ute
,
efter
som
de
nogsamt
kunde
finna
och
se
,
att
han
var
drucken
.

Lars
Mattsson
,
att
han
ingen
vidare
kundskap
har
om
Ekeroths
sjukdom
,
än
att
när
hans
hustru
i
veckan
före
påsk
var
hos
honom
och
han
frågade
efter
Ekeroth
,
skall
hon
svarat
,
det
han
1igger
sjuk
,
men
en
14
dagar
före
helgen
skall
han
varit
där
och
klagat
sig
över
en
stark
bröst
och
huvudsjuka
,
som
han
då
sade
sig
vara
besvärad
av
.

Responsum
,
av
skolmästaren
Brodenii
hustru
.

Qusestio
,
om
denna
Ekeroth
förr
pliktat
,
för
det
han
varit
drucken
?

Oansett
det
väl
kunnat
hända
,
att
denna
föravskedade
soldat
Erich
Ekeroth
haft
någon
känning
av
frossan
under
ottesångspredikan
nästlidna
påskdag
,
efter
som
han
förut
i
våras
varit
av
bemälde
sjukdom
besvärad
,
så
att
det
kunnat
föranlåta
honom
till
att
,
medelst
en
sup
brännvin
,
förekomma
sjukdomens
vidare
anfall
,
dock
emedan
han
intet
klagat
sig
för
någon
däröver
och
det
fördenskull
fast
likare
är
,
att
han
av
sin
efter
nämndens
intygande
vanliga
begärlighet
till
att
dricka
och
supa
gått
till
Hofgårdzberg
och
köpt
sig
brännvin
samt
supit
så
mycket
därav
,
att
han
blivit
drucken
,
var
med
han
så
mycket
mera
hade
bort
,
särdeles
emellan
predikningarna
på
en
så
stor
högtidsdag
,
innehålla
,
som
han
visste
,
att
han
intet
tål
stort
,
det
ock
,
när
han
fann
sig
så
beskaffad
,
hade
varit
bättre
,
att
han
hållit
sig
från
kyrkan
den
gången
,
än
att
han
skulle
gå
dit
och
göra
förargelse
;
Ty
prövar
tingsrätten
,
i
följe
av
Kungl.
Maij:tts
nådigaste
förordningar
om
svalg
och
dryckenskap
av
år
1733
och
dess
3
§
samt
om
oljud
och
förargelse
i
kyrkorna
av
år
1686
,
skäligt
,
det
bör
han
icke
allenast
,
för
det
han
varit
drucken
,
böta
sina
5
daler
silvermynt
eller
sitta
en
söndag
i
stocken
,
utan
och
,
för
det
han
kommit
drucken
i
kyrkan
under
gudstjänsten
och
gjort
förargelse
,
böta
sina
50
daler
silvermynt
eller
i
brist
av
bot
plikta
med
3
gånger
gatulopp
eller
,
så
framt
det
intet
bekvämligen
ske
kan
,
med
20
par
spö
till
3
slag
av
vart
par
samt
sedan
stå
uppenbara
kyrkoplikt
,
vilket
allt
dock
likväl
den
höglovlige
Kungl.
Maij:tts
och
riksens
Swea
Hovrätts
högtupplysta
och
nådrättvisa
omprövande
och
ändliga
utslag
i
all
ödmjukhet
underställt
var
/
Till
följe
av
vad
som
uti
förra
protokollet
finns
anfört
,
blev
den
grav
på
stora
gången
i
Wändels
kyrka
herr
häradshövdingen
Valtinsson
tillhanda
uppbjuden
andra
gången
,
som
han
köpt
av
postmästaren
Höök
uti
Yfre
för
sextio
daler
kopparmynt
.

Avskrivet
till
Kungliga
Hov
rätten
.

