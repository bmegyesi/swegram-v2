Blev
av
rätten
avsagt
,
det
en
syn
och
rådgång
nu
nästkommande
vårdag
hållas
skall
,
emellan
länsman
Måns
Andersson
i
Ede
på
den
ena
sidan
,
och
Sven
Olufsson
ibidem
på
den
andra
.

Anbelangande
intresse
må
söka
dem
i
Sundsvall
som
hans
gods
ifrån
honom
tog
.

(
19
)
Avsades
att
emedan
som
Erik
Nilsson
i
Näset
aldrig
har
köpslagit
med
Lars
Anderson
i
Rossiöö
(
?
)
om
alghuden
;
utan
med
hans
lagsmän
och
därför
dem
tillställt
6½
Rd:r
,
ty
kändes
han
fri
Larss
tilltalan
;
och
Larss
Andhersson
sökte
sina
lagsmän
som
huden
utom
hans
vetskap
sålt
ha
,
det
bäst
han
kan
och
gitter
.

Denne
Torkiel
har
icke
länge
varit
här
i
Jemptelandz
lappmark
,
utan
haft
sitt
tillhåll
uti
Ångermanlandz
lappfjäll
.

Var
uppå
strax
sjungs
Fader
vår
som
i
Himlen
är
/
eller
någon
annan
Psalm
;
Sedan
predikas
/
och
slutes
med
Bön
och
Välsignelse
.

Den
som
igenom
denna
större
Bannlysnlng
/
var
satt
utom
Guds
Församlings
gemenskap
/
skall
och
vara
utesluten
ifrån
alla
Samkväm
/
och
umgänge
med
annat
Folk
/
förutan
sin
Hustrus
/
Barns
och
Tjänstehjons
.

När
den
brottsliga
delen
/
som
för
Hor
/
ifrån
sin
äkta
Maka
skiljas
/
må
tillåtas
sig
att
gifta
/
och
med
vem
.
8
.

Vid
Äktenskaps
skillnader
/
brukas
följande
Formulär
:

Evangelium
eller
Lasten
,
som
efter
sedvänjan
plägar
i
Mässorna
lästa
eller
sjungen
vara
,
skall
man
ju
alltid
predika
,
så
väl
om
andra
Helgdagar
,
som
Söndagarna
,
och
ingens
helge
mans
Legendo
,
såsom
under
Påven
alltid
har
varit
sed
,
Ty
man
har
icke
många
sådana
Legendor
som
är
vissa
,
och
alldeles
komma
över
ens
med
Skrifterna
.

Dock
är
lika
mycket
vad
dessa
är
antingen
flera
eller
färre
,
män
eller
kvinnor
.

Så
förmanar
jag
,
att
man
för
all
ting
har
böner
,
åkallan
,
förböner
och
tacksägelse
,
för
alla
människor
,
för
Konungar
och
all
Överhet
etc.
Och
det
man
allramest
betänka
skall
,
så
har
ock
vår
HERre
Jesus
Christus
själv
satt
ett
dråpliga
stort
nådalöfte
till
den
allmänneliga
bönen
och
sagt
som
S
.
Mattheus
skriver
,
Där
två
av
er
komma
över
ens
på
jorden
,
vad
ting
det
helst
kan
vara
som
de
bedja
om
,
då
skall
det
dem
vederfaras
av
min
Fader
som
är
i
himmelen
.

För
all
mans
vittnesbörd
skull
,
och
till
att
förekomma
tvist
och
trätor
,
som
eljest
ofta
plägar
uppkomma
i
fästningar
,
skall
allmänt
ingen
fästning
ske
,
utan
in
för
Kyrkodörrarna
eller
i
Sakristian
.

Förfrågade
välaktig
Linnert
Jörensson
sig
här
för
rätta
om
Öckna
gård
,
således
att
all
den
stund
han
vänligen
var
förenat
med
Mats
i
Strengnäs
,
som
för
där
på
bott
hade
,
och
Lennart
undan
flydde
,
sedan
han
hade
sig
gården
avsagt
,
med
sådana
förord
,
att
när
Lennart
ville
flytta
från
gården
skulle
han
för:ne
Matz
samma
gård
hem
bjuda
,
vilket
och
med
skäl
och
bevis
skett
är
.

Kom
för
rätta
Hemingh
i
Båckabergh
och
Jon
i
Flahult
,
kyrkovärdar
i
Kårsberga
,
och
utfästa
samtliga
en
12
månne
ed
,
att
de
icke
till
det
ringaste
hade
för
snillat
av
Kronans
tionde
,
som
höge
överheten
welb:
Jöns
Larsson
till
Salzhult
hade
förlänt
.

Därmed
vart
han
för
båda
lägersmålen
sakfälld
till
penningar
—
60
marker
till
treskiftes
.

Då
med
vänlig
föraning
på
guds
och
överhetens
nådige
behag
med
härads
fogdens
,
nämndens
och
häradsmäns
samläggning
,
förlikades
Oluff
Karssonn
,
som
nu
bor
på
samma
gård
Nässiö
,
med
Jonn
Pärssonns
hustru
,
nämligen
Jngebor
Ericks
dotter
,
som
där
är
rätt
börd
till
jämte
vid
all
denna
släkt
,
att
han
för
nöjer
dem
alla
med
en
gått
vilja
12
daler
,
och
de
där
med
för
födda
och
ofödda
i
släkten
tillstå
och
tingsköta
honom
gården
efter
överhetens
nådiga
till
låtelse
att
bli
under
skatt
,
som
den
till
förne
warradt
har
.

Sakfälldes
Erich
Persson
Herr
Michilss
dräng
i
Börstill
till
—
3
daler
för
lytet
när
han
slog
sin
Matfaders
tänder
ut
fram
utur
Mun
,
och
till
—
20
₥
för
Shåremålet
:

Där
till
hustru
Margaretha
svarade
och
ville
bli
vid
sin
mans
Bok
,
och
alltså
skall
skulden
bli
mindre
.

kom
för
Rätten
Olof
Jönsson
ifrån
Norr
Tällghe
,
hustru
Charinss
ibidem
fullmäktig
,
och
gav
tillkänna
hennes
Man
Erich
Larsson
på
Singöön
död
bliven
vara
,
och
något
tillförende
kommen
i
Parlamentet
med
sin
halvbroder
en
borgare
ibidem
Michill
Jönsson
,
som
nu
flyktig
är
;
och
när
slagsmålet
skedde
bekom
hennes
Man
allenast
en
Pust
,
vilket
hon
föregiver
intet
vara
dödshugget
;
och
alltså
står
intet
på
sin
rätt
utan
vill
taga
förlikning
,
utan
annan
hastig
Sjukdom
skall
sig
sedan
ha
tillslagit
,
och
så
hårt
att
han
kom
ifrån
sitt
förnuft
förre
än
han
avsomnade
,
efter
som
Herr
Madz
Saccellanus
i
Häfröö
betygade
,
ty
för
hans
ursinnighet
skull
,
kunde
han
intet
med
dela
honom
Sakramentet
:

Johannis
tid
blev
han
igenhämtad
:
flera
vittnen
ville
Nillss
Persson
framha
men
nu
syntes
vara
Nog
.

Såsom
Hemming
Simonsson
i
Ränswed
,
har
lagt
en
Piga
Kerstin
Persdotter
från
Olof
Hindersson
i
Hohlborgen
förliden
Pingst
tid
,
skall
därför
plikta
3
mk:r
Sm:t
.
efter
15
Kap.
bygg:b
.
varmed
han
denne
gången
förskonas
.

Och
emedan
av
Nämnden
uppå
sin
eds
plikt
betygas
,
det
Finnäs
Hemmanet
är
kärandernas
rätta
börds
Jord
,
och
uti
deras
omyndige
år
,
är
dem
för
medelst
StugFaderns
vållande
ifrånkommit
;
Varför
erkänner
Rätten
skäligt
,
att
arvingarna
tillträda
Finnäs
hemmanet
igen
okvald
att
åtnjuta
för
sin
rätta
egendom
,
sina
utlagda
32
RD:r
igen
.

Till
detta
nekar
änkan
alldeles
,
sådana
ord
ej
ha
sagt
,
och
ej
heller
tillägger
änkan
Anders
vara
någon
baneman
Utan
sig
så
beklagat
,
att
Anders
var
hos
sig
samma
dag
och
velat
panta
sig
.

Enhälleligen
intygades
att
inga
oskattlagda
Allmänningar
här
i
Tinglaget
är
:
varandes
alla
avradsland
med
Rå
och
Rör
lagda
som
Specificerade
är
uti
Gamla
Böxlebreven
som
Anno
1666
dem
ifrån
tagna
blev
.

Anno
1729
den
29
September
,
hölls
efter
8
dagars
förutgången
pålysning
,
allmän
Mickelsmässo
Sockenstämma
,
med
St.
Malms
Församling
,
närvarande
Församlingens
Höge
och
Välborne
herrskaps
betjänter
,
Kyrkovärdar
,
Sexmän
och
meniga
man
,
då
efterföljande
av
slutat
blev
.
i
1
.

Och
emedan
,
sedan
Specialen
uppläst
var
,
på
de
fattigas
influtna
matvaror
,
många
fanns
,
som
aldrig
vilja
till
de
fattiga
förskjuta
,
besynnerligen
uti
Kåhlmårdz
Rootan
,
så
blev
de
närvarande
av
dem
,
allvarsamt
tilltalade
,
och
de
villiga
berömda
.
§
2
.

Icke
eller
vid
den
därpå
presenterade
och
igenomlästa
Specialen
på
FattigKassan
,
utan
befanns
alltsammans
ha
sin
riktighet
.

J
.
Dalenius
P
.
L
.
Nils
Nilsson
i
Bylen
Nämndeman
Pehr
Pehrsson
i
Stenta
Pehr
Pehrsson
i
Prästorp
Nils
Nilsson
i
Foglöö
Anders
Ersson
i
Foglöö
Jon
Swensson
i
Wråå

Och
som
Församlingen
ville
att
med
ett
nytt
taks
påläggande
,
fördröjas
skulle
till
vidare
,
blev
avslutat
,
att
de
gamla
bräder
skulle
i
höst
allenast
samman
jämkas
och
fastspikas
till
väggarnas
görligaste
konservation
.

Ehuru
allmänna
Sädesbristen
tycktes
,
å
ena
sidan
göra
saken
omöjlig
;
betraktade
likväl
,
å
andra
sidan
,
Församlingen
verkets
nödvändighet
,
och
i
anledning
därav
beviljade
,
att
taket
på
Tiondeboden
skulle
äntligen
bli
i
sommar
reparerat
,
och
så
mycket
av
den
fördärvade
ringmuren
omkring
Kyrkogården
,
som
förrådet
av
materialer
vill
tillsäga
$
16
.

Beklagade
Herr
Kyrkoherden
sig
,
mycket
,
att
avlidne
Soldaten
Kreymans
änka
hustru
Anna
,
ej
går
i
Kyrkan
,
samt
i
sitt
uppförande
på
ett
ohämmat
sätt
,
sig
oanständigt
skickar
,
utan
att
akta
de
enskilda
förmaningar
hon
titt
och
ofta
fått
.

Sven
Svensson
i
Karstorp
sexman
152

Gav
Herr
Probsten
vid
handen
,
att
utsocknesBor
på
sidstlidne
)
Vintertid
kört
in
med
sina
hästar
och
slädar
på
kyrkogården
bredvid
Magasins
huset
där
kyrkobalken
blev
riven
omkull
,
när
bemälda
Magasins
hus
uppsattes
;
Begärande
församlingens
tillstånd
att
få
,
med
den
grusen
som
tagen
är
utur
kyrkogården
till
gravlinjernas
hållande
,
låta
denna
öppning
på
KyrkoBalken
igen
täppa
och
mura
,
och
till
taket
därpå
betjäna
sig
av
den
spån
,
som
för
kyrkan
ligger
övrig
uti
MaterialBoden
,
vartill
församlingen
fann
sig
befogad
att
samtycka
.
§
9
.

På
träget
anhållande
,
beviljades
till
den
sjuklige
drängen
,
Eric
Jönsson
uti
Fiskartorp
,
12
dr
kmt
av
FattigKassan
,
till
underhåll
på
resan
åt
Medewi
Surbrun
,
under
lika
förbehåll
och
villkor
,
som
uti
förlidet
år
skedde
,
och
ses
pagina
)
304
.
§
15
.

Härpå
framkallades
både
Pehr
Jönsson
och
hans
Broder
Nils
i
Stensjö
,
såsom
ock
ovannämnda
drängar
,
och
frågades
Nils
,
vad
han
hört
av
Anders
Andersson
?

Att
så
tillgått
betygar
Fredrik
Tiselius
Gerhard
Lind
Pehr
Diuhlstedt
Pehr
Pehrsson
i
Brenäs
Olof
Pärsson
i
Benninge
Nämndeman
Kyrkovärd
Eric
Andersson
i
Mogetorp
Sexman

Och
kommer
denna
ordning
att
taga
sin
början
nästa
nattvardsgång
.
§
9
.

Vart
beslutat
och
av
gjort
,
att
Prästerna
vid
husförhören
skola
på
ett
särskilt
papper
noga
anteckna
alla
de
barn
,
som
innan
10:de
året
icke
lärt
läsa
rent
och
väl
i
bok
och
åtminstone
Luth.
Katekes
utantill
,
samt
att
dessa
barns
föräldrar
som
så
vårdslöst
barnens
uppfostran
,
skola
efter
en
och
annan
varning
plikta
2
dr
smt
,
vart
år
,
till
dess
barnen
lärt
sig
läsa
,
enligt
Kungl.
resolut
,
av
år
1723
.
§
6
.

Räkningen
upplästes
,
och
begärdes
pgr
därför
med
första
.

Stenqvists
hustru
,
som
lärt
2
gossar
i
Tiblenäs
,
att
läsa
i
ok
,
24
s.
S:a
22
R
.
40
s.
In
fidem
protokoll
Carl
F
.
Maneck
Den
14
juni
,
justerat
,
uppläst
,
erkänt
och
underskrivet
A
.
Lindblad

Augusti
)
1792
,
hade
denna
församlings
fattigkassa
tillfallit
105
R
.
36
s
(
sk
)
,
vilka
pgr
(
penningar
)
nu
å
kassans
vägnar
av
Prosten
emottogs
,
som
ock
kvitto
därpå
till
välbemälda
Herre
nu
överlämnades
.
3o
.

Ingrid
i
Mostugan
)
;
åbons
svärmor
i
Skräptorp
;
blinde
mannen
i
Nybygget
;
ä
.

Ingen
sockenhantverkare
begärde
avsked
.
§
6
.

Sålunda
vara
skett
,
intyga
å
församlingens
vägnar
undertecknade
Jac
.

Denna
lärdomen
om
Tron
,
var
hos
Aposteln
Paulum
allestädes
lärt
och
förkunnat
,
Såsom
till
de
Ephes
:
uti
det
2
Kap:
står
:

BEkännelsen
är
icke
heller
i
Guds
Församling
avlagd
.

I
förtiden
kom
de
tillsammans
i
Kloster
,
på
det
de
något
gott
skulle
lära
:

Borgmästare
och
Rådmän
för
sig
och
hela
Menigheten
.

Var
ofta
klagat
av
Stockholms
stad
/
Calmarna
/
Suderkoping
och
andra
Köpstäder
att
olaglig
köpslagning
sker
i
landet
/
städerna
till
fördärv
och
emot
lagen
/
då
man
vill
det
straffa
och
rätta
efter
lagen
/
falla
somliga
landsända
där
emot
och
vilja
att
sådant
icke
straffas
skall
/
och
följer
då
där
utav
/
att
om
man
i
de
måtte
gör
efter
lagen
/
skall
man
vänta
sig
uppstånd
och
obestånd
/
därför
gör
man
och
icke
efter
lagen
och
straffar
slika
oköp
bli
då
städerna
fördärvade
/
och
hela
landet
får
stort
oköp
/
och
vänds
dock
allt
Herren
till
/
att
han
det
vill
.

Detta
är
Riksens
Råds
brev
på
Westerårs
Recess
.

Till
att
bota
den
fjärde
bristen
/
samtycker
vi
alla
att
h
.
N
.
låter
bägge
parterna
av
lärarna
tillhopa
komma
och
disputera
i
vår
närvaro
/
att
man
måtte
höra
/
vilken
parten
rättast
hade
/
vilket
och
så
skedde
/
så
efter
vi
icke
annat
förnummit
antingen
av
samme
disputation
eller
av
deras
predikan
än
att
de
hade
god
skäl
/
och
icke
annat
predikade
än
Guds
ord
;
lovade
vi
h
.
N
/
att
med
det
rop
som
i
det
ärende
var
uppkommit
i
Riket
emot
h
.
N
.
var
i
sin
stad
stilla
ville
/
och
hjälpa
till
att
straffa
dem
som
sådant
falskeligen
utförde
Och
bad
där
alla
om
/
att
Guds
ord
måtte
allestädes
i
Riket
renliga
predikat
vara
.

I
Skolstugor
läses
efter
denna
Dag
Evangelium
ibland
andra
Läxor
/
efter
det
är
ju
Kristliga
Skolor
.

Lovade
taga
till
akta
.

Konung
Jahan
,
det
han
då
intet
eller
bevisa
kunde
vart
sagt
att
medan
den
Änka
där
boendes
är
kan
därför
göra
utlagorna
och
han
icke
visste
bevisa
sig
någon
bättre
rätt
där
till
skulle
hon
besitta
.

Anders
Andersson
Hock
Länsman
kärade
till
Per
i
Trosberga
om
5
t:nor
Säd
och
5
daler
9
T
/
s
öre
Penningar
,
vart
sagt
att
han
med
förste
skulle
betala
,
det
han
och
med
handslag
lovade
.

Vilken
hans
billiga
fordran
och
ingen
av
dem
för
vägra
visste
eller
kunde
,
och
fördenskull
enhälligen
vittnade
och
bekände
,
att
han
sig
där
sammastädes
,
såsom
en
Ärlig
Uppriktig
och
rättsinnig
man
ägnar
och
bör
väl
förhållit
hade
,
för
vilket
de
och
hade
orsak
honom
tacka
och
berömma
.

Dagsverken
nekade
Brundin
'
Åiwen
väl
till
och
sade
,
att
han
aldrig
förbundit
sig
där
till
.

Och
som
herr
kyrkoherden
i
följe
härav
anhöll
om
första
uppbudet
å
detta
hemman
i
Grytby
,
så
kunde
det
honom
intet
förvägras
,
efter
som
intet
klander
där
emot
förspordes
,
utan
blev
det
/
fördenskull
herr
kyrkoherden
tillhanda
uppbjudit
första
gången
.

Sedan
man
alltså
hade
hört
,
vad
han
härvid
kunde
ha
att
påminna
,
stannade
rätten
därvid
för
sin
del
,
att
bemälda
gästgiveri
,
som
består
av
ett
mantal
,
bör
och
kan
till
de
resandes
fortkomst
på
varje
fjärdedel
hålla
3
hästar
,
en
vagn
,
2
kärror
,
2
sadlar
och
2
slädar
samt
att
farten
intet
är
större
eller
trägnare
på
denna
vägen
,
än
att
bemälda
gästgiveri
väl
kan
vara
hållhästar
förutan
,
när
de
ha
och
hålla
så
många
hästar
i
beredskap
,
allenast
de
,
när
flera
erfordras
,
må
få
taga
hjälp
av
de
näst
omkring
liggande
byars
hästar
både
i
Norunda
och
Wendell
proportionaliter
,
samt
att
gästgivarna
,
som
är
tre
stycken
,
nämligen
Ohsengius
på
1
/
4
del
,
Lars
Jönsson
på
1
/
2
mantal
och
Erick
Jonsson
på
1
/
4
del
,
stå
varannan
bi
med
sina
hästar
,
som
de
efter
denna
nämndens
mening
kunna
hålla
,
vilket
ock
finns
vara
så
mycket
skäligare
,
som
de
alla
tre
formera
ett
gästgiveri
och
en
gästgivargård
.

Orkade
intet
bota
,
ty
avstraffades
hon
för
bemälde
40
daler
med
10
par
ris
till
3
slag
av
paret
40
Bonden
Oloff
Larsson
i
Kläringe
böter
,
för
det
han
utan
någon
orsak
eller
laga
förfall
absenterat
sig
ifrån
gudstjänsten
nästlidne
store
bönedagen
,
sina
10
daler
silvermynt
,
tilltalad
därom
av
Ikndzmannen
Gabriel
Wretberg
3
"
>
*
/
•
3
3
Unga
drängen
Erick
Persson
och
kvinnopersonen
Kierstin
Persdotter
i
Norrby
komma
för
otidigt
sänglag
med
varannan
att
erlägga
till
Wändels
kyrka
var
sina
2
daler
silvermynt
4
Mattz
Larsson
och
Anders
Erson
i
SkarpEkeby
är
sakfällda
,
den
förra
till
8
öre
och
den
senare
till
24
öre
silvermynt
,
för
förövad
olovlig
'
nävertäkt
uti
öhrby
frälse
säteris
hästhage
,
varom
de
blivit
instämda
och
tilltalade
av
befallningsmannen
Philip
Befvert
10V
.

