Länsmannen
Hans
Eriksson
Blix
anklagade
Faste
Larsson
i
Solberg
,
det
han
utom
laga
dom
har
inflyttat
sin
humblegårds
hage
in
på
sin
grannes
Sal
.

Efter
nämnden
av
de
12
saken
angick
,
remitteras
ärendet
under
landsens
24:s
dom
.

Angav
Jon
Nilsson
Ede
,
att
Olof
Svensson
i
Skerråsen
uti
olaglig
tid
,
emot
Kungl:
May:ttz
ordinantie
uppsåt
sina
älgs
led
,
dock
icke
honom
befunnit
någon
älg
att
ha
fått
.

På
bem:te
2:ne
års
ordinarie
räntor
till
6½
rd:r
8
sk:r
för
vartdera
året
,
vara
av
Måns
i
Moo
riktigt
betalade
och
kvitterade
på
befallningsmannen
sal
.

Så
emedan
Walle
och
Risselåhs
byägare
här
ifrån
sig
ej
undandraga
kunna
,
så
vara
till
gånget
;
utan
för
Rätten
,
tillika
med
tolvmän
tillstå
och
bekänna
så
uti
fordom
dagar
varit
;
men
förmedhelst
manfall
på
be:te
Joenssgården
,
är
det
så
ej
uti
akt
tagit
dessutan
draga
så
väl
Jonss
Gårdsman
lika
skatt
till
Kungl:
May:tz
och
kronan
,
efter
sina
tundl:d
,
med
all
där
av
gående
besvär
och
tunga
,
som
östbyggare
Walle
och
Risselåhs
män
för
sina
tundl:d
.

Men
hans
börda
och
mössa
fanns
strax
igen
i
sjön
ett
stycke
ifrån
byn
,
och
igen
liknelse
till
själva
personen
.

Befinnes
ett
extrakt
av
Hammerdahls
kyrkoböcker
avkopierat
och
vidimerat
av
lagman
sal
.

Olof
Abrahamsson
som
okallad
lade
sig
uti
en
annans
sak
och
förde
osanning
att
Jon
Sjulsson
ej
var
stämd
,
som
dock
övertygades
av
länsman
och
Jöns
Eriksson
i
Sikås
vara
stämd
,
sakfälldes
till
3
m:k
Sm:tt
efter
29
kap.
kungs.b.ll
.

Oluf
Siulsson
föregiver
vara
här
till
lockad
och
övertalad
av
fältvebeln
Lars
Hindriksson
,
då
han
reste
till
Norrige
,
som
fick
honom
2
dukater
och
2
Rd:r
med
det
förord
,
om
han
skulle
få
tobaken
i
Norrige
på
kredit
,
skulle
han
ha
hem
penningarna
6
Rd:r
vilket
Oluf
Siulsson
i
god
trohet
gjort
och
visade
honom
sina
specie
penningar
,
då
Lars
Hindrichsson
där
emot
upptog
6
Rd:r
i
karoliner
att
ombyta
,
fick
således
fält
vebeln
sina
penningar
igen
.

Kyrkoherdens
hustru
beklagar
sig
och
bortmist
2
klimpar
smör
som
hon
saknar
vilka
konan
Anna
Olufzd:r
har
stulit
och
det
inlagt
uti
sin
systers
Sara
Olufzd:rs
kista
,
om
söndagen
medan
folket
var
i
kyrkan
har
hon
in
krupit
genom
fönstret
,
och
det
uttagit
och
lovat
till
sockenstuge
hustru
,
Brita
Larsdotter
,
vilket
smör
beräknas
till
1
(
pund
)
har
de
alla
3
bytt
sin
emellan
som
värderas
till
1:16
öre
.

Erik
Månsson
i
Fyrås
har
genom
länsman
i
Lit
stämt
Hemming
Sjulsson
i
Ytter
Näset
för
det
han
har
förhållit
pigan
Kerstin
Wellamsdotter
gå
i
tjänsten
,
men
ej
kommit
tillstädes
,
sakfälldes
efter
33
kap.
ting
b
LL
3
m:kr
.

Löjtnanten
utvalde
Erik
Samuelsson
,
Daniel
Andersson
och
Jon
Olofsson
i
Hallen
.

Om
allmänningarna
rannsakades
och
befanns
att
fyra
st.
finnar
har
sig
nedersatt
inemot
Ångermanlandz
gränsen
och
1680
blev
de
skattlagda
och
rörlagda
och
flera
boställen
finnas
och
där
sammastädes
.

Jon
Olofsson
i
Gåxsjö
angav
hurusom
han
på
Daniel
Olofssons
hemman
ib:m
fått
för
14
à
15
år
sedan
dom
brev
,
vilket
2
à
3
år
därefter
medelst
en
skadlig
vådeld
uppbrann
och
ty
begär
att
han
må
kunna
sig
till
säkerhet
få
å
nyo
ett
dombrev
,
vilket
Daniel
Olsson
tillstår
och
ånyo
köpsedel
givit
och
många
kunnigt
;
ty
skall
i
protokollen
där
efter
rannsakas
och
likmätigt
det
11
kap.
Jordb
.

Soldaten
Mathias
Dreflingh
och
Bärent
Musicant
hjälpte
honom
dricka
ur
ölkannan
och
efter
honom
blev
och
sig
lade
kvar
.

Soldaten
Mattias
Jacobsson
Åbergh
skuldgavs
ha
belägrat
Märit
Persdotter
ifrån
Goxsjö
som
födde
barn
förliden
Larsmässo
.

Anna
Mårtensdotter
i
Öhn
hans
där
insatte
3½
kanna
brännvin
i
h
.
Vellams
hustrus
namn
uttagit
och
uppdruckit
,
det
Nills
tillstår
och
säger
sig
vara
förlikt
därom
och
skall
giva
på
sin
part
3
d
.

Såsom
Ramsehlerne
föregiva
sig
efter
Olof
Persson
och
Ingemar
Erikssons
i
Vallen
och
Erik
Zakrissons
i
Tärsjö
begäran
allenast
dem
till
skogs
följt
och
ej
kunna
annat
förstå
än
att
de
pretenderade
2ne
älgsdjur
fälldes
inom
Ångermanlandz
landamäre
och
Giörwijkerne
påstå
det
vara
skett
inom
Jemptelandz
landsskrå
,
varför
kan
intet
slut
däruti
ske
,
förr
än
orten
och
hullstan
blir
i
ögnasyn
tagna
,
var
av
prövas
kan
på
vars
skog
djuren
fällda
är
och
ty
lämnat
till
syn
och
besiktning
.

Var
till
med
är
Nills
Ståckman
som
förvites
med
hust
.

Allt
så
kan
Rätten
för
denna
gången
saken
icke
slutligen
avhjälpa
utan
till
nästa
laga
ting
uppskjuta
,
då
Nills
Swartt
skall
förpliktat
vara
sina
vittnen
i
saken
ha
tillstädes
och
dom
avvakta
.

Drar
och
någon
hit
in
Lärare
av
en
främmande
Religion
,
till
någon
Gudstjänsts
övning
/
eller
till
Barns
undervisning
i
Religionen
;
så
skall
den
samme
böta
/
till
nästa
Hospital
eller
Husarme
500.de
Dahl:r
Silvermynt
/
och
förvisas
Riket
.

Såsom
en
noga
Uppsyn
med
Ungdomens
upptuktelse
/
Studier
och
Resor
i
främmande
Land
/
drar
i
längden
efter
sig
en
stor
nytta
/
för
Guds
Församling
och
det
världsliga
Regementet
/
och
lätteligen
hända
kan
/
medan
de
vistas
ibland
Folk
av
villfarande
Religioner
,
att
de
och
insuga
villfarande
Meningar
/
dem
de
sedan
oförsiktigt
bringa
med
sig
hem
i
Landet
igen
/
sig
och
andra
till
skada
och
fördärv
;
Alltså
förmanar
Vi
alla
/
i
synnerhet
Föräldrar
/
eller
dem
som
stå
i
Föräldrars
stad
/
och
vilja
sända
sina
Söner
eller
Förvanter
i
främmande
Land
så
och
dem
själva
/
som
är
komna
till
sina
myndiga
år
/
och
av
eget
Råd
/
vilja
sig
en
slik
Resa
företaga
/
att
först
och
främst
bära
åhåga
om
det
/
som
till
deras
Själs
Salighet
länder
/
vinnlägga
sig
om
vår
Kristliga
Religions
rätta
Kunskap
och
övning
/
och
vad
som
där
till
hör
/
samt
noga
underrätta
sig
/
om
ovanberörda
Slut
och
Stadgar
/
på
det
de
så
mycket
bättre
må
veta
att
vakta
sig
för
främmande
Gudstjänster
/
hålla
sig
stadigt
vid
Guds
heliga
Ord
/
och
undfly
deras
umgänge
/
som
söka
att
bedraga
dem
ifrån
vår
rätta
/
till
någon
villfarande
Lära
.

§
.
I
.
Prästerna
skola
flitigt
/
fram
för
andra
/
läsa
den
heliga
Skrift
/
och
troligen
bedja
Gud
/
om
Nåd
och
Upplysning
/
att
de
den
samma
må
rätteligen
kunna
förstå
/
och
så
tiIl
sin
egen
/
som
sina
åhörares
Bättring
och
Salighet
/
lära
och
förklara
.

Prästen
blottar
allenast
Barnets
Huvud
/
och
det
med
Vatten
begjuter
/
brukandes
där
vid
de
Ceremonier
och
Böner
/
samt
det
sättet
/
som
här
till
dags
varit
vanligt
/
och
uti
Handboken
infört
är
.

Vill
Syndaren
/
av
fruktan
för
Straffet
/
sig
där
till
intet
bekväma
/
och
Synden
är
av
den
Art
och
Natur
/
att
hon
är
fullbordad
/
och
intet
mer
kan
lända
till
någons
fördärv
och
skada
/
då
skall
Predikanten
något
dröja
med
avlösningen
och
Herrens
Nattvard
/
med
mindre
Syndaren
är
stadd
i
Dödsfara
:

§
.
I
.
Ehuruväl
Vi
våra
Undersåtar
/
emot
allehanda
Missgärningar
/
Laster
och
Odygder
/
med
god
Lag
/
Ordningar
och
Stadgar
/
således
försett
har
/
att
den
Processen
,
som
till
Bannlysning
hör
/
med
den
högstes
Bistånd
/
ej
någon
tid
/
eller
fast
sällan
/
skall
behövas
;
Likväl
/
såsom
det
i
första
Kristliga
Kyrkan
har
varit
brukligt
/
så
är
och
nödigt
/
att
vid
någon
sådan
händelse
/
i
vårt
Rike
/
Guds
Kyrka
och
Församling
/
vilkens
uppsikt
/
vård
och
försvar
/
av
Gud
oss
anförtrott
är
/
må
veta
/
hur
där
med
skall
förhållas
/
är
om
Bann
således
stadgat
/
som
följer
.

Avstår
han
ändå
intet
med
Synden
/
då
må
omsider
hans
Kyrkoherde
/
sedan
Sakens
sannfärdiga
beskaffenhet
/
är
oss
först
och
förut
vorden
kungjord
/
och
han
/
uppå
Biskopens
och
Konsistoriets
befallning
/
har
/
tre
Söndagar
i
rad
/
lyst
honom
till
bättring
/
upptäckt
hans
fel
/
och
förmanat
Församlingen
/
att
bedja
Gud
för
honom
/
alldeles
avsöndra
en
så
förhärdad
och
obotfärdig
Syndare
/
ifrån
Guds
Församlings
gemenskap
/
och
uppenbarligen
av
Predlkstolen
Bannlysa
honom
/
på
efterföljande
sätt
:

Men
när
så
fordras
/
att
någon
ny
Bön
skall
författas
/
och
till
en
viss
Tid
brukas
/
då
bör
Ärkebiskopen
/
tillika
med
Consistorio
Ecclesiastico
,
efter
Vår
Befallning
/
henne
på
ren
Svenska
/
med
Gudliga
Ord
/
förutan
Prål
och
vidlyftiga
Omsvep
/
sammansätta
/
och
Oss
tillhanda
sända
/
då
Vi
vill
den
samma
överse
låta
/
och
sedan
till
Stiften
skicka
/
att
brukas
i
Församlingarna
.

Om
någon
Tvist
uppkommer
/
vilken
rätta
Giftoman
är
/
eller
och
den
samme
missbrukar
sin
Makt
och
Myndighet
.
3
.

När
Tvist
blir
om
själva
Trolovningen
/
samt
Gåvorna
.
4
.

När
skillnad
sker
i
Äktenskapet
/
vem
som
bör
förse
de
Barn
/
som
bägge
Föräldrarna
kännas
vid
/
och
vad
vars
och
ens
Giftorätt
är
/
uti
boet
som
skall
skiftas
.

Men
likväl
må
Parterna
dem
i
DomKapitlen
först
angiva
/
och
där
försökas
/
om
en
god
och
vänlig
förlikning
kan
ingås
/
uti
de
mål
/
som
kunna
och
böra
förlikas
.

Giftermål
med
främmande
Religions
Förvanter
/
måste
flitigt
avrådas
;
Dock
blir
de
icke
alldeles
förbjudna
/
för
Hoppet
om
deras
omvändelse
/
till
Vår
lära
/
och
när
de
ingås
med
sådana
villkor
/
som
Våra
Stadgar
påbjuda
.

Men
om
det
ej
vinnas
kan
/
hänvisas
de
till
världslig
Rätt
/
där
att
rannsakas
och
dömas
om
själva
Gärningen
/
var
utur
skälet
till
skillnaden
sökes
.

§
.
V
.
Om
någon
efter
Trolovningen
/
egenvilligt
reser
ifrån
sin
Fästmö
/
och
emot
hennes
samtycke
/
blir
länge
borta
/
må
henne
tillåtas
/
att
gifta
sig
med
en
annan
;
Dock
skall
hon
först
giva
sig
an
hos
Biskopen
och
Konsistorium
.

När
en
eller
två
blir
besmittade
uti
ett
Hus
/
då
skola
de
andra
strax
Gudeligen
och
väl
bereda
sig
/
till
att
begå
HErrens
Nattvard
/
tillika
med
den
Sjuka
.

Nyfödda
Barn
/
som
icke
har
satt
Döpelsen
/
för
deras
hastigt
avgång
skull
/
skola
njuta
deras
Föräldrars
Lägerstad
/
och
Prästen
vara
där
tillstädes
/
tiIl
att
kasta
Mull
på
dem
/
och
läsa
en
Bön
.

Förgriper
sig
någon
här
emot
/
så
skall
han
därför
tillbörligen
ansedd
bli
och
plikta
.

Om
Valet
faller
på
någon
som
icke
är
dess
värdigare
/
och
Biskopen
finner
/
att
i
Stiftet
andra
är
/
som
de
intet
känna
/
vilka
för
sin
lärdom
/
långliga
Tjänst
/
goda
Gåvor
och
Skicklighet
/
böra
fram
för
den
de
åstunda
/
med
befordran
ihågkommas
/
de
där
gott
Vittnesbörd
om
sig
ha
/
och
giva
det
säkra
hoppet
/
att
Församlingen
igenom
dem
skall
märkligen
kunna
uppbyggas
och
förkovras
;
Då
böra
de
i
det
som
skäligt
är
/
och
till
deras
bästa
länder
/
låta
rätta
sig
/
och
åtnöjas
med
Biskopens
och
Konsistoriets
Förordning
Försummar
någon
Församling
/
i
rättan
tid
/
denna
sin
nödtorft
för
Biskopen
att
andraga
/
så
måste
han
/
uppå
Prostens
härom
gjorde
påminnelse
/
utse
för
dem
en
tjänlig
/
god
och
trogen
Kyrkoherde
/
tagandes
med
sina
Kapitels
Män
för
sig
anteckningen
på
de
äldste
/
lärdaste
och
bäst
förtjänade
Skolbetjänter
/
Krigspräster
/
och
Kapellaner
i
Stiftet
/
som
vänta
efter
laglig
Kallelse
till
bättre
Lägenhet
/
och
där
av
föreslå
en
eller
två
/
som
bekvämligast
prövas
/
det
lediga
Rummet
att
förträda
/
dem
de
dit
förskicka
/
att
göra
prov
Predikan
/
och
inhämta
Församlingens
samtycke
och
ordentliga
Kallelse
;
var
uppå
sedan
StadfästelseBrev
av
Biskopen
skall
meddelas
.

Men
om
Valet
är
fallet
på
en
värdig
Man
/
emot
vilken
Biskopen
ej
har
sådant
Jäv
som
sagt
är
/
då
bör
han
sätta
honom
till
den
föreslagna
Lägenheten
.

Men
här
till
höra
då
alla
ordningar
,
som
gå
på
vissa
och
bestämda
tider
och
bekvämlig
rum
,
när
och
varest
Kristet
folk
sig
församla
skall
,
då
allmänneligt
Predikan
,
Böner
,
Sakramenten
,
och
vad
annat
sådant
är
för
Kristligt
handel
,
Ty
efter
detta
icke
allestädes
kan
ske
var
dag
,
eller
uti
all
rum
,
kräver
nöden
här
med
en
viss
ordning
,
sådana
som
varit
har
,
icke
under
Påven
allenast
,
utan
ock
eljest
i
hela
Kristenheten
,
med
beskedda
dagar
,
dem
man
nu
nämner
Helgedagar
.

Item
,
Att
allt
det
som
i
Församlingarna
handlas
,
skalvtrettas
på
allmänt
förståndliga
mål
.

Och
har
den
meningen
varit
hos
alla
Kyrkornas
Lärofäder
,
att
sådana
besvärjelser
skall
vara
kraftigt
emot
djävulen
.

Efter
vilkas
goda
och
Kristliga
exempel
ock
så
några
Gudfruktiga
Svenska
Konungar
sig
tagit
har
,
läggandes
sig
där
mycket
ut
om
,
att
Kristen
tro
ock
så
här
i
Swerige
skulle
planterat
och
utspridd
varda
,
Såsom
nämligen
den
förste
Konung
Biörn
,
vilken
genom
inkallade
Predikare
S
.
Ånsgarium
och
andra
,
här
i
Riket
lät
predika
Kristen
tro
.

Så
är
ock
icke
heller
det
nyttigt
,
att
de
enfaldiga
sig
bekymra
med
mångahanda
Postillor
,
som
nu
nog
är
förhanden
,
och
dagliga
mer
förökas
,
Ty
där
med
varda
de
mer
förbistrade
och
hindrade
,
än
till
det
de
mena
,
förfordrade
,
och
förlöper
än
då
dess
förinnan
tiden
,
vilken
de
eljest
till
att
själva
begrunda
och
överväga
saken
,
Ja
ock
till
att
läsa
något
tjänligt
stycke
i
Skrifterna
,
med
stor
fördel
bruka
måtte
,
Ty
är
ock
måttan
här
uti
god
,
så
att
man
råder
sig
en
Postillo
den
som
rättsinnig
är
,
eller
åt
mest
två
,
och
låter
sig
där
med
nöja
,
och
brukar
Skrifterna
desto
bättre
.

Item
,
Där
utinnan
är
min
Fader
prisat
,
att
ni
bär
mycket
frukt
.

Efter
som
ock
i
Psalmen
står
,
Gud
säger
till
den
ogudaktiga
,
Hur
förkunnar
du
mina
rätter
etc.
Ty
ligger
ock
då
största
makten
där
uppå
,
att
Predikarna
själva
frukta
Gud
,
vilket
om
de
rättsliga
göra
,
varder
han
dem
givandes
,
både
det
,
att
de
visliga
tala
(
såsom
han
lovade
Aposteln
,
sägandes
,
Jag
skall
giva
er
mun
och
visdom
etc.
Och
att
med
deras
tal
följer
lycka
och
salighet
.
,
,
,
,

Item
ock
så
(
det
långt
för
vår
tid
av
kommet
var
)
honung
,
mjölk
.

Så
behålla
och
bruka
Kristna
församlingar
än
nu
för
samma
sak
skull
några
av
dessa
gamla
Ceremonier
,
sommestädes
flera
och
sommestädes
färre
,
efter
som
väl
möjlighet
är
att
ske
må
,
först
man
denna
deras
grund
vet
,
och
ger
icke
dem
mer
tillförne
än
det
sig
bör
,
eller
håller
dem
så
enkom
vara
av
nöden
,
såsom
meningen
under
Påvens
regemente
varit
har
och
än
nu
hos
de
enfaldiga
mycket
vara
gitter
,
varför
ock
Prästerna
skola
här
om
fliteligen
undervisa
meniga
man
,
att
de
slika
tankar
här
om
icke
ha
skola
,
Eljest
lika
som
en
part
av
dessa
Ceremonier
hos
oss
för
denna
saken
skull
är
bortlagda
,
så
kan
det
samma
ock
väl
ske
med
flera
där
av
,
där
man
icke
vill
låta
sig
här
om
rätt
undervisa
.

Men
givs
ock
sådana
svar
,
att
man
icke
kan
vara
fullviss
uppå
om
barnet
är
rätt
döpt
eller
ej
,
Då
skall
det
icke
dess
heller
döpas
under
villkor
,
såsom
de
Påvska
icke
rätt
lärt
och
gjort
har
,
sägandes
,
Astu
icke
döpt
,
så
döper
jag
dig
etc.
Ty
sådana
dop
har
ingen
rätt
och
Kristlig
art
,
utan
man
skall
uti
sådana
fall
döpa
villkorslöst
,
alldeles
såsom
man
eljest
plägar
,
och
Döpelsens
rätta
grund
kräver
.

Till
det
andra
hör
vi
här
ock
,
vad
både
barnen
och
vi
har
för
en
stor
tröst
,
nämligen
,
att
Guds
Son
Jesus
Christus
vår
Herre
så
redebogen
är
till
att
hjälpa
alla
dem
som
till
honom
komma
,
vare
sig
ung
eller
gammal
,
Så
att
han
ock
storliga
tog
dem
till
vedervilja
som
slikt
med
denna
barnen
förhindra
och
icke
tillstädja
ville
.

Sedan
de
har
rättat
sig
upp
igen
,
frågar
han
barnens
namn
,
och
tar
så
vatten
i
händena
,
och
gjuter
tre
resor
över
barnens
huvud
,
sägandes
.

Och
där
han
av
alla
dessa
befinner
att
barnet
är
rätt
döpt
,
skall
han
låta
bli
där
vid
,
och
ingalunda
döpt
på
nytt
,
Ty
det
är
ett
Dop
och
icke
flera
,
såsom
S
.
Paulus
betygar
,
Utan
han
skall
sådana
Dop
gilla
,
och
uti
allas
deras
åhöro
som
då
är
tillstädes
,
stadfästa
med
slik
ord
som
här
efterfölja
.

Efter
det
första
slaget
,
skriftade
sig
Publikanen
i
Templet
,
och
eljest
otaliga
många
flera
,
som
Skriften
omtalar
,
Vilka
alla
ock
där
igenom
fullkomliga
fått
har
syndernas
förlåtelse
,
Ty
är
hon
ock
lika
som
av
Gud
befallet
,
rätteliga
av
nöden
,
så
att
henne
förutan
kan
platt
ingen
komma
till
syndernas
förlåtelse
.

Dock
var
dess
förinnan
några
av
dem
något
förekommer
,
som
Pastor
loci
behöver
veta
.
det
skall
han
honom
kungöra
.

Var
några
framkomma
till
Skrift
,
som
så
är
till
ålders
komna
,
att
dem
bör
veta
och
kunna
läsa
Fader
vår
,
Tron
,
Bodhorden
etc.
och
han
som
Skriftemålen
hör
,
befinner
att
de
slikt
än
nu
intet
kunna
,
Då
skall
han
desto
flitigare
förmana
dem
,
att
de
sådant
än
nu
med
det
allraförsta
lära
,
så
att
de
ock
ingalunda
bjuda
sig
fram
till
Sakramentet
,
för
än
de
det
allt
redliga
har
lärt
och
kunna
.

Sedan
skall
man
ock
fråga
honom
till
som
Skriftemålen
gör
,
om
han
begär
varda
avlöst
.

Men
efter
det
till
åtskillig
brott
hör
ock
åtskillig
plikt
,
Ja
,
ock
väl
till
åtskilliga
personer
i
samma
sak
,
hör
åtskillig
plikt
,
kan
icke
väl
någon
allmännelig
form
eller
sätt
här
uppå
givet
warda
,
Ty
måste
det
ock
mest
stå
till
hans
förnuft
,
beskedlighet
och
trohet
,
som
Skrifterna
sätter
.

Kristliga
Sekvenser
må
man
ock
undertiden
sjunga
,
särdeles
på
dessa
högtider
,
Jul
,
Påsk
,
Helge
Torsdag
och
Pingstdag
.

O
Barmhärtige
himmelska
Fader
,
uti
vilkens
händer
står
allt
världsligt
våld
och
överhet
etc.
Men
efter
detta
sättet
är
uti
så
måtto
endel
för
långt
,
när
man
har
Messan
för
händer
,
är
det
avkortat
,
och
brukas
nu
allmänt
så
,
att
man
vart
stycket
strax
efter
det
andra
uppräknar
sägandes
.

Till
det
nionde
begär
Rauall
,
att
det
måtte
rannsakas
,
hur
otroligen
Linnert
handlade
med
99
års
skaffuell
fläsk
,
som
samme
år
borde
utgöras
,
och
prövas
vad
kronan
där
av
bekommit
har
,
ty
där
som
det
hade
blivit
levererat
till
Calmare
,
måtte
räkenskapen
det
utvisa
.

På
samma
sätt
förmäler
Rauall
,
att
han
har
handlat
med
en
bonde
i
Alzeda
socken
,
benämnd
Anders
i
Ödshult
,
vilken
Anno
98
gav
Linnert
ena
ko
i
mjugg
,
så
släpade
han
med
två
oxar
till
kronan
,
för
det
hans
hustru
hade
haft
lägersmål
och
gjort
hor
med
en
dräng
,
Sunderbo
Nils
benämnt
.

Vad
Godskalcks
gods
anbelangar
,
som
Linnert
Jörensson
skulle
vederkänts
efter
för:ne
Godskalck
Jonsson
,
som
uttrymde
,
om
vilket
Raffuall
begär
fullkomlig
veta
besked
,
vart
allt
sådant
var
tagit
vägen
.

Och
på
denne
försäkring
förtalade
bonden
för
sin
själa
herde
,
huruledes
han
hade
sett
en
gräslig
gärning
,
som
ganska
ohövligt
var
till
att
omtala
.

Men
någon
tid
där
efter
begynte
åter
prästen
samme
handel
innerligt
att
begrunda
och
revolvera
huruledes
han
sig
här
utinnan
skulle
rådföra
,
alldenstund
för:nB
hans
socken
bonde
,
som
honom
sådan
handel
i
tromål
hade
uppenbarat
,
var
en
sanningsman
,
där
för
måste
och
hans
ord
och
tal
följa
skäl
.

Och
där
på
gav
han
mig
fyra
skilling
etc.
Till
vilket
drängen
alldeles
nekade
att
han
dem
skamlig
gärning
icke
hade
bedrivit
.

Samma
dag
begärde
en
av
nämnderna
,
Hans
Håkonsson
i
Tälleridh
här
för
rätta
av
häradshövdingen
och
nämnden
,
att
hans
jord
;
brev
på
Tällerids
gård
och
dess
torp
stad
måtte
varda
renoverat
och
förnyat
,
vilket
jorda
brev
Michill
Sigfridson
hade
utgivit
Anm
1571
Uppbudna
Gårdar
Allan
västra
gården
i
Byestadh
i
Alzeda
socken
30
Allan
Brunns
gården
i
Bexeda
socken
2
°
Allan
Göliarids
gården
i
Korsberga
socken
2
°
Allan
östra
Endagarden
i
Nye
socken
2
°
Allan
Ödzhulte
gården
i
Alzeda
socken
2
°
Allan
västra
gården
Trälarp
i
Nyjo
socken
2
°
Allan
gården
Mösshult
i
Alzeda
socken
1
°
Allan
gården
Hesleåsa
i
Stenebergh
socken
i
°
En
hel
sättnings
gård
i
Högakull
i
Alzeda
s.
2
°
1
/
2
gård
i
Endarydh
i
Byrcke
socken
1
°
1J2
gård
i
Endarydh
i
Alzeda
socken
2
°
En
hel
gård
Störriarp
i
Stenebergh
socken
i
°
En
frälse
gård
Lambåsa
i
Alzeda
socken
30
En
skatte
utgjord
i
Faderstårp
i
Nye
socken
30
ANNO
CHRISTI
1602
den
11
augusti
stod
laga
härads
ting
Österherrat
å
rätta
tingstad
uti
närvaro
ärlig
och
välbördig
]
Jöns
Larssons
till
Salzhult
,
välförståndig
Linnert
Jörenssons
i
Hunde
stad
,
kronans
befallningsman
i
för:110
härad
,
välaktig
Suen
Månsson
i
Rösa
underfogdes
samt
hederlige
och
vällärde
mans
här
Gudmund
i
Kårsberga
.

Kom
för
rätta
en
knekt
hustru
,
benämnt
Sigridh
i
Måshult
i
Rampnkulla
socken
och
klagade
på
Nils
i
Bexeda
,
att
han
hade
släppt
en
tjuv
olagvunnen
,
som
hade
henne
ifrån
stulit
svart
blaggarn
19
alnar
.
vadmal
13
alnar
,
ringare
ett
kvarter
,
penningar
2
Va
nw£er
,
sundeskt
en
aln
,
vantar
3
par
,
ett
ärmekläde
och
några
band
.

Men
efter
hon
inlät
sig
med
honom
till
en
vänlig
förening
Edemän
hans
.

Emellertid
kom
grevinnans
gods
fogde
dit
,
som
han
sig
sedan
inflyttat
hade
,
och
ville
utkräva
återstädjan
och
veta
för
vad
orsak
han
var
olagligen
med
åminne
av
flytt
hennes
gods
.

Men
var
han
icke
allt
som
föreskrivet
står
efter
hans
tillsägelse
och
förpliktelse
efterkommer
och
fullbordar
,
skall
hans
dom
och
straff
stå
honom
öppen
före
.

Kom
för
rätta
Måns
Jngesson
i
Boda
,
och
klageligen
gav
till
känna
,
att
hans
granne
Anders
Jutte
ibidem
icke
ville
bli
vid
den
förlikning
dem
emellan
lagligen
med
bägges
deras
vilja
och
samtycke
gjort
var
;
och
vite
var
dem
emellan
satt
,
att
vilken
förlikningen
först
avbröt
,
skulle
böta
3
oxar
och
3
daler
,
och
nu
bevisades
att
Anders
Jutte
hade
avbrutit
,
och
för:ne
Måns
hårdligt
till
livet
undsagt
,
evar
han
honom
överkomma
kunde
,
och
vart
därmed
till
vitet
fälld
.

Brynell
i
Nyaby
i
Alzeda
socken
fullmyndig
på
Oluffs
vägnar
i
Häsleåker
och
på
alla
Oluffs
syskons
vägnar
,
nämligen
Gummes
i
Broby
i
Laneskeda
socken
,
Jngridis
och
Jngebors
vägnar
i
Näffuelsiö
och
på
Marrietes
vägnar
i
Diuranäs
i
Byrke
socken
,
så
och
fullmyndig
på
Bengt
Nilssons
vägnar
i
Näsiö
i
Huetlanda
socken
,
så
och
fullmyndig
på
Oluff
Carlssons
hustru
vägnar
ibidem
,
Elines
nämligen
,
och
på
Segrid
Nilsdotters
vägnar
ibidem
.

Och
var
Jon
Persson
i
Såndåker
fullmyndig
på
Oluff
Lassessons
vägnar
i
Gältarid
i
Myresiö
socken
,
på
Segrid
Lassesdatters
vägnar
ibidem
och
på
Jngrid
Lasses
dottors
vägnar
i
Brantas
i
Näffuelsiö
socken
.

Därmed
avhänder
han
nu
ifrån
sig
och
sina
arvingar
för:ne
halva
Store
Ödzhulte
gård
,
och
till
ägnar
den
in
under
Suen
Månsson
hans
barn
och
rätte
efterkommande
arvingar
etc.
Kom
för
rätta
Nils
Jonsson
i
i
Slätåkra
i
Alzeda
socken
fullmyndig
på
sin
hustrus
Bengtas
vägnar
,
så
och
fullmyndig
på
Håkones
vägnar
i
Trijshilt
i
Myresiö
socken
och
på
Suens
vägnar
i
Såndåker
i
Bexeda
socken
,
att
tingsköta
Jöns
Sigfridsson
i
Endegården
i
Myresboda
i
Nya
socken
Jöns
Erickssons
,
Oluff
Erickssons
och
Jngofredes
del
i
för:ne
gård
,
som
är
en
treding
av
halvan
för:ne
gård
,
för
et
par
oxar
,
ena
ko
,
en
fyra
lod
silver
sked
och
penningar
efter
deras
eget
goda
nöje
för
rätta
köpt
,
och
sex
mark
i
ettleffue
för
samma
treding
.

Kom
för
rätta
Per
Matsson
i
Snuggarp
i
Skyre
socken
samt
Per
Halffuarsson
ibidem
med
deras
hustrur
,
barn
och
allt
sitt
husfolk
och
var
i
synnerhet
gjorde
sin
ed
på
lagboken
att
de
aldrig
vetat
,
hört
eller
sett
hade
någon
liknelse
eller
besked
till
,
att
Per
Matsson
i
Snuggarp
,
skulle
ha
burit
hem
,
eller
förnummit
att
han
,
eller
någon
i
hans
hus
något
rådjur
skulle
ha
förtärt
,
sålt
eller
bort
gömt
,
som
Håkon
Månsson
i
Loaklöff
föregivit
och
berättat
har
.

Och
samma
natt
kom
hon
sin
kos
.

Men
alldenstund
Rauall
icke
till
det
ringaste
i
samma
sina
beskyllningar
kunde
med
vittne
eller
skäl
Linnert
Jörensson
överbetyga
,
att
han
någon
otrohet
eller
orättrådighet
H:F:N
.
eller
kronan
hade
bevisat
,
utan
nämnden
och
menige
häradsmän
med
uppräckta
händer
gav
honom
ett
uppriktigt
och
ärligt
skottsmål
,
att
han
troligen
och
rättrådligen
,
både
emot
högbe:lt
höge
överheten
och
eljest
emot
var
man
här
i
häradet
i
sin
tillbetrodde
befallning
sig
skickat
och
ställt
hade
.

Kronans
befallningsman
välbemälde
Linnert
Jörensson
uppbjöd
sig
i
menige
mans
åhöro
och
närvaro
,
om
någon
här
i
häradet
fanns
,
som
honom
vad
som
helst
skänk
eller
gåva
hade
givit
eller
förärat
och
till
det
ringaste
där
över
hade
till
att
kvida
,
då
ville
han
den
,
nu
i
sin
välmakt
,
samma
skänk
efter
likmätig
värdering
okvidande
igen
vederlägga
.

Kronans
befallningsman
ärlig
och
välförståndig
Linnert
Jörensson
uppbjöd
sig
efter
samma
sätt
som
på
tinget
näst
tillförne
.

Varför
tillsporde
herr
Erich
Peer
Ravaldzson
i
Elmesta
,
varför
han
det
talet
har
utkommit
där
till
han
Nekade
,
men
herr
Erich
beropade
sig
på
en
Student
benämnd
Andreas
Gåse
,
som
skall
om
detta
vara
hans
sagesman
,
där
till
Per
Ravalsson
nekade
,
därhos
var
bemälde
Andreas
intet
tillstädes
,
därför
blev
Saken
uppskjuten
:
vad
Säden
anlangar
som
för
herr
Erich
bortkom
,
bekände
han
sig
den
eljest
ha
utur
släden
förtappat
,
och
gjorde
bemälde
Olof
fri
,
men
om
utslagna
öga
skall
vidare
rannsakas
.

Då
svarade
bemälde
herr
Madz
att
bemälde
Anderss
tog
två
tunnor
Råg
av
honom
för
10
år
sedan
,
då
galt
tunnan
10
daler
Nu
begärde
Anderss
tillstånd
att
leverera
honom
Säd
igen
;
men
Herr
Madz
svor
högeligen
sig
ha
honom
Säden
levererat
för
betalningen
.
där
till
Anderss
Nekade
,
ej
heller
fanns
vittne
där
till
:
varför
avdömdes
,
att
herr
Madz
skall
betala
Anderss
Jönsson
sina
penningar
,
igen
uti
sådant
mynt
som
han
det
tog
,
eller
annat
vitt
Mynt
efter
Riks
Daler
värde
;
när
bemälde
gäll
gjordes
,
och
Anderss
betalade
åter
herr
Mattz
,
Rågen
i
penningar
,
för
så
myket
herr
Matz
skäligen
bevisa
kan
tunnan
gullit
ha
enär
den
gällen
gjordes
,
medan
Anderss
intet
bevisa
kan
sig
ha
allenast
tillsagt
honom
Säd
igen
och
intet
penningar
61
.

Orsaken
till
käromålet
är
att
enär
bemälde
Salig
Olof
tjänade
för
bemälde
hemmanet
Sättra
,
högg
han
på
deras
Skog
Svedjeland
,
där
förbrände
han
några
Ekar
;
därför
fordrar
välborne
Jonas
Bureus
böterna
av
Sättraborna
;
Varför
förmenade
Madz
Madzson
sig
ville
igen
något
vinna
av
hans
arv
;
Där
till
bemälde
Per
i
Bredhsättra
svarade
,
sig
mera
gäll
för
sin
bemälde
broder
betalat
ha
,
än
det
värt
var
som
fanns
efter
honom
;
Och
medan
bemälde
Oloff
för
Riksens
fiender
på
platsen
bliven
är
,
skall
här
om
först
bevis
givas
till
Höge
Överhetens
vidare
förklaring
.
66
.

framkom
Peer
i
Stridzby
,
och
anklagade
Olof
i
Lervijken
,
som
efter
sin
Sons
döds
avfall
hade
hans
lösören
borttagit
,
och
intet
sin
bemälda
Sonhustru
,
som
är
bemälde
Perss
dotter
därav
antvardat
.
som
var
ett
åketyg
,
2
pund
Lin
,
och
några
penningar
.

Där
till
Nekar
han
alldeles
att
han
gör
Kamstadh
by
något
intrång
på
Mulbeethen
,
medan
torpet
där
han
nu
är
,
ligger
fjärran
där
ifrån
.
7
.
vad
den
lille
Ängen
anbelangar
som
nu
bärgas
till
Torpet
,
sade
han
sig
vilja
bruka
bönen
och
söka
om
han
henne
åtnjuta
kunde
.
8
Föregiver
han
sig
ha
Salig
Mårthen
Jacobssonss
tillstånd
att
bygga
på
Kamstadh
ägor
sedan
han
själva
hemmanet
avträdde
,
därpå
han
intet
skriftligt
uppvisa
kunde
,
utan
beropade
sig
på
välaktat
Engellbrecht
Svänsson
och
Thomass
i
Myrby
uti
Danmarks
Socken
uti
vilkas
Närvaro
,
han
skall
honom
det
ha
tillstått
,
varför
blev
här
med
dilaterat
till
dess
skriftligt
besked
ifrån
dem
uppvisas
.
85
.

Och
alldenstund
hon
ingen
skrivelse
ifrån
honom
bekommit
har
,
var
hon
sinnat
till
att
inlåta
sig
uti
Äktenskapet
med
bemälde
Madz
Persson
Och
medan
hon
intet
Lagligen
eller
vidare
förra
än
hon
lät
sig
belägra
,
har
efterfrågat
om
sin
mans
86
.
död
,
därhos
befanns
klarligen
av
de
besked
som
Abraham
Olofzson
,
krigs
Cammarerer
och
Anderss
Persson
Humble
,
utur
Rullarna
som
i
den
höga
Kungl.
Krigsrätt
finnas
utgivit
ha
,
den
ena
daterad
29
december
1636
,
och
den
andra
7
April
Anni
huius
,
vilka
klarligen
utvisa
att
bemälde
hennes
man
har
levat
,
och
var
då
under
välborne
herr
Åkee
Hanssons
etc
Regemente
,
Varför
dömdes
bemälda
Anna
och
Matz
Persson
ifrån
livet
,
efter
Guds
Lag
,
Genesis
6
.
etc.
Dock
dess
Höglovlige
K
.
Hovrätts
förklaring
förbehållen
.

blev
efter
dess
höglovlige
Kunglige
hovrätts
förklaring
,
utgiven
13
oktober
1634
av
Nyio
rannsakat
om
det
dråpet
som
Johan
Mårthensson
i
Rissby
uti
Vixsta
Socken
,
en
Ryttare
,
på
en
annan
Ryttare
benämnd
Peer
Haansson
i
Ahlbärgha
uti
Vändel
Socken
begått
har
,
sedan
denne
Peer
hugg
fått
hade
,
fördes
han
till
bemälde
Rissby
,
Låg
där
till
Sängs
i
fyra
dygn
,
gick
uppe
sålänge
som
här
efter
förmäles
,
brände
sig
själv
i
ett
sår
med
ett
glödhett
Järn
,
att
en
åder
mera
uppkom
,
och
därför
begynte
blodet
mera
än
tillförne
rinna
;
vilket
ärende
är
till
Vändels
Ting
remitterat
,
till
att
där
av
Nyio
rannsakas
,
dock
där
intet
upptagit
,
alldenstund
Peer
Haansson
sig
här
uti
Häredet
bränt
har
,
där
och
eftertecknade
vittnen
boendes
är
:
vilka
åtskiljeligen
förhördes
,
och
efter
Eds
å
bok
avläggande
således
vittnade
som
följer
:

När
han
så
länge
som
bemält
är
till
Sängs
legat
hade
,
och
till
att
Läkas
antagen
av
Johanss
Svärfader
Olof
Hollm
,
gick
han
mestadels
uppe
in
till
bemälde
tid
Då
Johanss
Bröllop
hållit
blev
,
där
han
ibland
andra
gjorde
sig
lustig
.

När
hon
bemälde
brände
sår
jämte
de
andra
förbundit
/
:
hon
var
och
understundom
där
tillförne
men
intet
då
han
brände
sig
:
/
begynte
blodet
att
stiga
uppföra
och
armen
svartna
varigenom
stor
värk
förorsakades
,
Per
bad
för
Guds
skull
att
hon
ville
lösa
upp
såret
som
förbränt
var
,
när
det
skedde
,
sprutade
blodet
såret
,
och
långt
ifrån
utan
någon
uppehållning
,
åter
förband
hon
det
,
strax
begynte
Per
Haansson
kvida
,
intill
dess
det
upplöstes
,
och
blodet
sedan
stadigt
rann
,
När
hon
det
sista
gången
om
Torsdagen
förbundit
hade
sade
han
,
löser
upp
det
det
blir
likväl
min
död
,
med
samma
förbindande
höll
hon
fort
fyra
gånger
om
dagen
.

Samma
dagen
,
uppsteg
för
Rätten
dess
Ädles
och
välborne
111
.

Anders
som
mest
i
Humbleö
uppfödd
var
,
kom
till
gården
-
S
.
Jacobj
tid
,
Då
Lovade
han
salig
herren
tiänst
,
icke
allenast
till
Mickels
mässo
,
utan
och
sedan
;
Olof
svarade
att
drängen
,
hade
intet
stått
sig
till
tjänst
.

Oloff
svarade
sig
intet
där
av
veta
,
En
tid
där
efter
kom
Oloff
Stille
ifrån
Staden
och
sände
bud
efter
Anderss
,
vilken
strax
begav
sig
ifrån
gården
till
honom
,
och
intet
tänkte
på
sitt
förra
Löfte
,
och
hade
sedan
mest
sitt
tillhåll
i
bemälde
Muthsunda
,
och
förde
ved
till
Stockholm
att
försäljas
,
En
tid
där
efter
blev
kunnigt
var
han
var
,
dock
vidare
intet
efter
honom
frågat
,
förra
än
den
18
.

S
.
dagen
framträdde
för
Rätten
hans
Nådes
herr
Päer
Baners
etc.
Fullmäktig
,
Mortenn
Hanssonn
,
och
kärade
till
Johann
i
Knuteby
Länssmann
,
om
någon
gälsgårds
till
ett
hundrade
famnar
som
han
hade
bortfört
,
ifrån
Långarnn
Äng
,
och
den
sig
till
nytta
avhänt
,
Där
till
Johann
svarade
,
att
medan
han
tillförne
hade
sin
målgård
kring
om
bemälde
Äng
,
ty
ängarna
vore
intet
ändå
åtskilda
,
Nu
har
han
samt
hans
grannar
dem
åtskilt
,
är
och
Tälge
Stad
intresserat
med
Knutebyess
äng
.

Varför
begärde
han
dilation
,
till
dess
de
opartiska
vittnen
som
över
Kontraktet
vore
komna
tillstädes
,
som
vetskap
här
om
ha
skola
,
Såsom
veta
betyga
om
Mäster
Bärendt
några
Penningar
på
handen
tagit
har
,
när
de
efter
avlagda
Ed
,
här
om
vittna
,
varder
Saken
vidare
som
vederbör
utförd
.
121
.

framkom
Engelbrecht
de
Vretz
och
själv
bekände
sig
ha
för
2
år
sedan
fört
på
sin
Skuta
åt
Dantzick
några
stänger
Fransos
Järn
,
dock
honom
oveterligen
,
till
vilket
han
föregav
sina
Båtsmän
Erich
Jonsson
,
Per
Månsson
och
Olof
Nillsson
svara
skola
,
och
det
för
Arrendatorerna
var
de
Järnet
bekommit
ha
.

Saken
av
vägen
:
vilka
klagomål
skola
i
lika
måtto
hans
Nåde
Landshövdingen
andragas
.

Såsom
hon
det
ville
avslå
:
/
sådant
intet
värt
vara
.

Varför
gav
de
sin
Kyrkoherde
Herr
Måånss
i
Löffsta
sådant
tillkänna
,
vilken
förmanade
dem
till
att
taga
förståndiga
kvinnor
,
som
henne
rannsaka
skulle
,
det
de
och
gjorde
,
sände
bud
efter
hustru
Dårdhi
i
Åkerby
och
hustru
Brijta
ibidem
dessa
vittnade
efter
eds
avläggande
,
sig
finna
sådana
Mjölk
uti
hennes
Bröst
,
Såsom
den
där
Nyligen
fött
hade
ha
Plägar
;
Därhos
var
hon
ändå
svullen
över
livet
,
vilket
de
sade
och
ett
visst
tecken
där
till
vara
.

När
hon
nu
som
bemält
är
för
Rätta
hades
,
stod
hon
i
förstone
på
sin
förra
bekännelse
,
och
ville
intet
ut
med
sanningen
,
ehuru
hon
där
till
med
flit
och
foglighet
förmanades
:
då
blev
och
henne
förhållit
vad
bemälda
kvinnor
hos
henne
rannsakat
och
funnit
hade
,
och
ytterligare
på
åtskilligt
sätt
förmanad
sanningen
bekänna
;
Då
svarade
hon
sig
bli
belägrat
av
bemälde
Anderss
S
.
Mickelsmässo
tiden
,
och
fått
missbörd
distings
tiden
,
som
sig
skall
förorsakat
ha
av
det
hon
lyfte
Säden
på
PörthessLaffuan
,
och
alldenstund
det
hade
ingen
Skapnad
,
kastade
hon
det
i
ugnen
:
än
förhölls
hon
på
sätt
som
förre
,
och
förmanades
till
sanningens
bekännelse
:

Och
kunde
intet
Rätten
för
detta
uti
Saken
till
dom
skrida
,
ej
heller
bemälde
Henrich
värja
eller
fälla
,
förra
än
de
tillstädes
komma
,
1
som
såg
när
gossen
hugg
fick
.
2
de
som
honom
sedan
synat
har
,
både
medan
han
levde
,
och
sedan
han
död
blev
.

Efter
långsamt
övervägande
Döms
Jöns
Larson
till
12
mk:r
efter
det
4
Kap:
i
S:M
:
med
våda
Blev
och
in
för
rätten
med
Handband
förlikt
att
Jöns
Larson
skulle
giva
Änkan
Anna
Edfwardzdotter
hustrun
till
den
döde
Otta
RD:r
.

Framkallades
vittnen
som
inne
var
,
när
dråpet
skedde
,
Erick
Gudmundson
och
Jöns
Gudmundson
i
Hemsiöö
,
berättade
att
Erick
Jonson
som
dräpt
blev
,
slog
Faltin
Jacobson
ett
munslag
och
sade
detta
skall
du
ha
för
Källar
nyckeln
;
Den
dräptes
Syster
Anna
Jonsdotter
,
bekände
ock
att
Sahl.Erick
Jonsson
sade
till
Faltin
,
detta
munslag
skall
du
ha
För
Källar
nyckeln
,
Och
vill
du
mera
ha
så
skall
du
få
,
och
med
det
samma
slog
han
honom
med
en
Kniv
i
hjärtat
,
och
följde
honom
,
fort
efter
in
åt
stugan
,
till
dess
han
sig
på
sätet
nedsatte
,
var
efter
han
och
strax
gav
upp
andan
.

Efter
denne
avsagde
dom
faller
Dråparen
Jöns
Pehrson
till
ödmjuk
bön
,
så
hos
gud
först
som
sedan
hos
den
höge
Överhet
om
nåd
och
lindring
på
straffet
,
helst
emedan
han
och
sig
med
den
döde
\
emellertid
som
han
levde
/
så
som
och
målsäganden
förlikt
har
,
att
han
sin
rätt
honom
godvilligt
tillgivit
har
som
är
att
se
av
\
ett
/
Kontrakt
\
som
de
sig
emellan
slutit
/
(
10
RD:r
)
\
har
,
och
han
det
ännu
in
för
rätten
tillstår
/
rätten
det
bekänner
,
att
han
intet
strävar
efter
hans
liv
för
sin
person
;
Utan
hemställer
det
alltsammans
den
höglovlige
Kungl:
Hovrätts
höga
betänkande
och
gunstiga
resolution
,
vad
straff
helst
\
den
/
sig
behagar
\
och
för
gott
finner
/
att
han
under
gå
måtte
.

Erick
Erickson
i
Finnäs
låter
uppbjuda
Wästergården
Flattnor
2
gången
.

Brodde
Olufsson
i
Anwijken
,
Oluff
Nilsson
i
Öbyn
,
Lars
Broddesson
i
Backe
,
Jon
Nilsson
i
Gåssböhle
Lars
Larsson
i
Bensiöö
,
Erich
Larsson
i
Anwijken
,
Erich
Pehrsson
i
Flatnohr
,
Jon
Pehrsson
i
Bossiöö
Pehr
Jönsson
vid
Ån
,
Nilss
Nilsson
i
Mordwijken
Mattes
Pehrsson
i
Fanbyn
och
Oluff
Andersson
i
Wärwijkn
.

Gästgivaren
i
Brek
Swän
Nilsson
Lät
uppbjuda
Salmon
Larssons
gård
i
Benssöö
halv
annan
tunnland
Jord
Ibidem
Andra
gången
.

Allmogen
\
i
Bräcke
/
begärde
Delation
av
Herr
Befallningsmannen
om
kärrorna
till
att
förfärdiga
till
våren
och
bli
alltså
förskonade
att
de
ej
mer
skulle
böta
än
var
man
3
mk:r
och
Gästgivare
6
mk
Sven
Nilsson
i
Bräcke
6
mk
Ty
där
finns
allt
odugliga
Kärror
så
att
den
vägfarande
Man
som
för
Penningar
Leja
vill
Lider
stort
och
män
och
bräck
Utlovandes
bot
och
bättring
.

(
42
.
)
Sammaledes
Peder
Bengtsson
i
Marsätt
och
Sundsiöö
Socken
,
Trädde
för
Rätten
,
(
uppbjudandes
½
Tunnland
i
Landsom
,
tredje
gången
för
40
RD:r
Köpt
)
Presenterandes
sin
sal
.

Besvärade
sig
vördige
Kyrkoherden
vällärde
H:r
Isaac
Alstadius
,
öf:r
sina
åhörare
i
Bräcke
Socken
,
undantagandes
gästgivaren
Swän
Nillsson
har
på
Kungl.
Kommissorial
rannsakningen
i
Rödhöön
hos
Richz
Rådens
Hög
wälb:ne
H:r
Gustaf
Posse
och
H:r
Johan
Gylldenstierna
utverkat
sig
på
orätt
berättelse
en
Resolution
att
de
skulle
föra
sin
korntionde
allenast
till
Bräcke
Kyrka
och
icke
på
Offne
,
där
för
kyrkobords
ägor
tillbytt
är
,
efter
Riks
Rådets
Högvälborne
H:r
Claes
Stiernskiöldz
nådgunstige
Disposition
,
att
bruka
kyrkobord
blev
bytt
till
Krono
Jord
där
gästgivaren
Swän
Nillsson
åbor
och
Kyrkoherden
bekom
Offne
i
stället
för
Bräcke
Kyrkobord
,
dit
de
är
pliktiga
föra
sin
Korn
tionde
,
dock
likväl
uti
anseende
så
Procederat
är
,
så
proponerade
vördige
kyrkoherden
att
Bräcke
bönderna
må
på
läggas
efter
Kungl.
Krögare
ordinatier
få
för
penningar
leja
deras
hästar
,
att
de
be:te
sin
tionde
må
föra
till
Offne
som
är
Bräcke
kyrkobord
vilket
vördige
Kyrkoherden
sådant
ej
kan
lagl
.
förvägras
,
utan
de
må
sig
där
efter
rätta
.

Tobaks
besökaren
Jonas
Pehrsson
,
angav
det
Joen
Olufsson
i
Grimnäs
har
handlat
med
Tobak
och
det
köpt
av
Oluf
Kopparslagares
son
,
Erich
där
av
sålt
Johan
Olufsson
par
alnar
,
och
när
han
skjutsade
besökaren
,
sålde
han
honom
½
aln
Såsom
dessa
sig
här
ifrån
ej
unddraga
kunna
Utan
tillstå
så
vara
tillgånget
,
Varför
efter
Maij:ttz
Plakats
12
.
punkt
sakfälldes
vartdera
...
8
D:r
Sm:tt
;
Men
Johan
Olufsson
äger
intet
att
böta
med
,
ty
skall
han
plikta
med
fängelse
.

Anders
Erichsson
i
Rijse
ifrån
Lockne
Socken
beklagade
sig
det
Oluf
Hansson
i
Böhle
har
för
någon
tid
sedan
beskyllt
honom
ha
mördat
och
ihjälslagit
Pehr
Persson
i
Hööwijken
ifrån
Båssiö
Socken
,
var
till
Oluf
Hansson
nekar
ej
så
ha
sina
ord
fällt
;
Länsman
Pehr
Anderss
vittnade
det
sal.Pehr
Persson
i
Hööwijken
har
för
4
år
sedan
1675
fört
Kyrko
tionden
till
Prästgården
har
han
varit
i
länsmansgården
då
han
var
Krankaktig
och
svullen
i
ögonen
av
den
sjukdom
nembl:n
Fransos
han
var
bekaiadt
med
,
då
begivit
sig
till
h
.
Sara
Prästänkan
i
Skoron
där
han
över
Natts
låg
,
och
morgonen
där
efter
,
kört
med
störste
eländighet
hem
\
ifrån
/
Skoron
,
som
var
1
mil
emellan
,
där
han
under
vägen
är
död
bliven
och
hästen
drog
honom
hem
på
Släden
till
sin
gård
.

Emot
Länsman
Pehr
Andersson
och
Pehr
Bengtssons
Söner
,
Angående
Sundz
Hemmanets
Inlösen
,
vilka
bägge
stämdes
till
nästa
Laga
ting
med
sina
brev
och
vittnen
.

B
förmäler
Ty
kunde
Rätten
Saken
ej
längre
uppskjuta
,
Utan
Länsman
Pehr
Andersson
har
efter
19
och
22
kap:
ting
b
.

Jöns
Jonsson
i
Ösiö
,
uppbjuder
halva
hemmanet
som
hans
broder
barn
tillkommer
,
första
gången
pantsatt
för
43
RD:r
2
.
20
.

Item
Inkaminerade
Pastor
en
Kopia
av
Kungl.
Maij:tz
Resolution
given
Prästerskapet
i
Jemptelandh
d
.
25
September
Anno
1668
och
dess
8:de
punkt
av
innehåll
att
de
Skogar
,
ängar
och
fisken
som
kunna
tillförne
antingen
av
Sueriges
eller
Dannemarckz
Konungar
och
Biskopar
Prästerskapet
Och
Kyrkorna
förunnade
vara
,
att
de
konserveras
och
förblir
vid
deras
rätta
ägare
med
nådig
vilja
att
Guvernören
,
Prästerskapet
i
den
provinsen
som
i
den
andra
allt
görligt
assistans
bevisar
,
havandes
och
Prästerskapet
Lag
och
Rätt
för
för
!
sig
uti
den
Landsorten
.

Och
alla
ingen
Särdeles
skatt
därför
göra
utan
hålla
före
,
att
skatten
på
deras
Hemman
är
förd
,
för
givandes
bem:te
Personer
det
hela
Fiällstadh
med
Råå
och
Röör
är
belagt
,
Oluff
Pärsson
berättade
det
Erich
Jonsson
efter
1646
års
dom
intet
bekom
Fiällstadh
,
utan
måste
lösa
sin
Svärfaders
Jöns
Gelofssons
Systers
Barbrus
Arvs
part
där
uti
,
Av
Peder
Jönsson
i
Torwalla
och
Brunflod
Socken
som
Barbrus
Dotter
till
hustru
bekom
.

Iag
skall
skrubba
er
för
än
denna
Aktion
ändas
,
och
att
han
intet
vill
eller
kunde
gå
in
medan
Fänriken
där
var
,
eftersom
han
hotades
med
sin
värja
göra
dråp
;
Fänriken
bekände
sig
allenast
säga
om
jag
icke
fick
ligga
där
inne
så
skulle
han
det
göra
Protesterandes
emot
Fänrikens
Förvitelse
i
sin
Inlago
,
görandes
bli
vid
Sveriges
lag
och
Präst
privilegierna
Maintinerat
.

Sist
förbjudes
och
dem
alla
till
fång
,
som
icke
till
Kvarn
byggningen
i
synnerhet
nödiga
är
att
röra
och
tillgripa
,
vid
laga
Plikt
tillgörande
.

Malmgryttan
föregiver
han
sig
köpt
av
Hust
:

Dito
,
och
omsider
utfästa
18
D
.
Sm:t
,
var
med
h
.
Kapten
lät
sig
benöja
,
och
Mickell
sträckte
Kapten
hand
där
över
,
att
betala
till
S
:

Och
ändå
dem
icke
borde
lidne
,
eller
efterlåtit
varda
,
sig
här
i
Riket
nedsätta
,
som
med
någon
falsk
Lärdom
umgå
,
och
med
oss
uti
Läran
icke
ens
är
,
på
det
de
andra
med
sig
icke
förföra
måtte
:

Sedan
igenkommandes
till
att
döma
levandes
och
döda
.

Vilken
för
oss
människor
,
och
för
våra
salighet
skull
,
nedersteg
av
himmelen
,
och
tog
mandom
genom
den
heliga
Anda
,
av
Jungfru
Maria
,
och
vart
en
människa
:

ITem
varder
lärt
,
att
det
är
en
helig
Församling
,
den
ock
alltid
bli
skall
.

ÄNdock
Guds
Församling
egentligen
är
de
Heligas
och
rätte
Kristtrognas
Samkväm
:

Sammaledes
förkastas
ock
de
som
lära
,
att
syndernas
förlåtelse
,
icke
givs
genom
tron
,
utan
bjuda
,
att
man
Guds
nåd
förtjäna
skall
genom
våra
egna
förnöjelser
.

Dock
förstör
icke
Evangelium
världsligt
Regemente
och
Hushåll
,
utan
alldeles
befaller
,
att
man
allt
sådant
hålla
och
bruka
skall
,
såsom
Guds
egen
ordning
,
och
uti
sådana
stånd
bevisa
den
Kristliga
kärleken
.

Därför
har
våra
Predikanter
,
om
Tron
,
Guds
Församling
således
lärt
och
undervisa
som
nu
följer
:

Varför
ock
Christus
säger
hos
Johannem
i
det
15
Kapit
:

Men
den
heliga
Skrift
lär
intet
att
vi
skola
tillbedja
eller
åkalla
framlidna
Helgon
,
eller
ock
av
framlidna
Helgon
hjälp
söka
och
begära
.

Men
det
har
varit
en
allmännelig
klagan
,
att
några
missbruk
skola
hänga
hos
gemena
Kyrkostadgar
:
varför
efter
dessa
missbruk
,
med
gott
samvete
icke
kunna
gillas
,
är
de
mestadels
förändrade
vordna
.

Det
samma
vittnar
ock
Hieronymus
,
vilken
säger
:

Varför
,
om
några
vilja
heller
annamma
bägge
delarna
i
Herrens
Nattvard
,
borde
dem
icke
varda
tvingadhe
att
de
annorlunda
måtte
göra
,
med
deras
samvets
besväring
.

Men
om
Mässan
utplånar
de
levandes
och
dödas
synder
,
för
det
omak
och
arbete
,
man
har
till
att
höra
henne
,
så
bekommer
man
rättfärdigheten
därför
,
att
Mässan
hålls
och
hörs
,
och
icke
igenom
Tron
,
vilket
den
heliga
Skrift
ingalunda
lida
kan
.

Men
denna
Pauli
lära
,
är
nästan
platt
utsläckt
vorden
av
människo
stadgar
,
vilka
har
denna
mening
av
sig
fött
,
att
man
igenom
åtskillnad
på
mat
,
och
andra
sådana
stadgar
,
ändliga
måtte
förvärva
nåd
och
rättfärdighet
.

Item
Paulus
till
de
Romare
i
det
14
Kapit
:
säger
:

Dock
likväl
behålls
hos
oss
mestadelen
av
de
stadgar
,
som
tjänliga
är
där
till
,
att
all
ting
mante
uti
Guds
Församling
skickligt
tillgå
:

Till
det
första
,
varder
hos
oss
lärt
,
att
det
är
alla
efterlåtit
giva
sig
i
Äktenskap
,
som
icke
bekvämliga
är
,
till
att
vara
det
förutan
,
för
ty
Klosterlöften
kunna
icke
förstöra
eller
omintet
göra
Guds
bud
och
ordning
.

Om
man
nu
detta
dem
till
förtret
ville
skärpa
och
driva
,
hur
mycket
kunna
man
finna
och
sammanhämta
,
där
själva
Munkarna
nu
skämmas
vid
?

OM
Bisparnas
kall
och
ämbetes
kraft
,
är
i
förtiden
mycket
vordet
disputerat
:

Vilket
de
tog
uti
beråd
och
på
sistone
fullo
till
och
både
honom
/
att
han
skulle
stå
fast
uti
det
som
han
då
företagit
hade
emot
K
.
etc.
Och
sade
h
.
N
.
till
hulskap
och
manskap
/
lovandes
vilja
stå
med
honom
med
liv
och
makt
/
så
efter
h
.
N
.
sagt
att
där
ingen
var
som
regementet
ville
taga
sig
före
/
och
farligt
var
att
icke
skulle
vordet
fullföljt
till
ändan
det
företaget
var
/
anammade
då
h
.
N
.
regementtet
i
Guds
namn
och
gjorde
där
om
så
mycket
honom
möjligt
var
och
efter
som
Gud
gav
nåden
till
.

Först
att
samme
ed
och
bepliktelse
har
h
.
N
.
av
somliga
intet
varit
hållen
utan
aldrig
snarare
Riket
var
kommet
i
sin
frihet
igen
/
begyntes
strax
stämplas
obestånd
och
förräderi
emot
h
.
N
.
där
han
dock
aldrig
med
hans
vit
någon
tillfälle
tillgivit
hade
/
som
var
först
med
Mäster
Knuth
och
h
.
Peder
Canceller
/
vilka
h
.
N
.
i
förstone
beslog
där
med
och
dock
såg
utöver
med
dem
för
goda
mäns
bön
skull
/
förhoppandes
att
de
skulle
bättra
sig
/
och
sedan
har
sådant
fördrag
/
som
de
och
satte
goda
män
i
borgen
för
sig
/
att
det
icke
mer
ske
skulle
/
vilket
de
dock
intet
hålla
/
utan
när
h
.
N
.
var
faren
till
Dannmarck
på
Riksens
bästa
/
att
förhandla
om
frid
och
endräkt
emellan
Riken
/
förgät
icke
samme
Mäster
Knuth
och
h
.
Pedher
deras
förräderi
/
utan
fullföljde
det
/
givandes
sig
upp
i
Dalarna
/
stämplandes
där
uppresning
emot
h
.
N
.
diktandes
på
honom
många
oredliga
stycken
som
breven
väl
utvisa
som
de
kring
om
landet
skrivna
/
efter
vilket
de
och
på
sistone
rättad
vorde
/
för
vilka
saker
h
.
N
.
satte
ett
allmänneligt
möte
här
i
Westeras
/
och
bevisade
här
för
den
meneman
slika
stycken
vara
honom
oredliga
pådiktat
och
ljugen
/
och
var
då
åter
redebogen
att
övergiva
regementet
att
för
h
.
N
.
skuld
icke
skulle
behövas
något
obestånd
företagas
i
Ritket
.

Ibland
annat
det
h
.
N
.
så
påförs
är
detta
ett
/
om
de
hjälper
som
förlidna
år
har
pålagda
varit
att
de
för
ofta
ske
/
den
ena
efter
den
andra
/
den
mene
man
till
fördärv
etc.
Det
bekänner
h
.
N
.
att
samme
hjälper
är
oftare
på
lagda
en
h
.
N
.
ville
/
för
den
feges
skuld
h
.
N
.
haft
har
sedan
han
kom
till
regementet
emot
K
.
etc.
Söffrin
Norby
och
andra
hans
parti
:

Sammalunda
ropas
och
om
Gripzholms
Kloster
att
h
.
N
.
det
nederlag
/
är
Er
mesteparten
väl
alla
vitterligt
att
det
var
och
är
h
.
N
.
arv
och
eget
/
och
vart
utan
hans
faders
vilja
emot
lagen
skickad
till
Kloster
/
och
är
klart
att
om
h
.
Sten
Sture
hade
haft
barn
/
hade
det
visserligen
aldrig
vordet
Kloster
/
därför
stod
h
.
N
.
väl
till
att
bygga
det
.

Item
:
var
det
icke
hjälpa
kan
/
förs
då
h
.
N
.
uppå
att
han
indrager
nya
tro
i
landet
/
det
dock
h
.
N
.
förstånd
har
/
att
Kyrkans
förmän
med
deras
anhang
honom
mest
pådiktad
ha
/
fördenskull
att
h
.
N
.
och
jämväl
många
andra
så
nu
här
som
i
flera
andra
Riken
har
lärt
befinna
många
stycke
där
Kronan
Riddarskapet
och
den
meneman
av
Kyrkans
personer
har
med
bedragna
och
förtungade
varit
/
vilka
med
tiden
väl
förtäljda
varda
/
och
har
med
slika
stycken
upphävt
sig
för
Herrar
underkuvad
landsens
Furstar
/
Riddarskapet
och
den
meneman
/
slagit
under
sig
samt
med
självdiktade
Gudstjänst
/
den
Gud
aldrig
bjudit
har
samt
pantat
köpet
överlåtit
.
etc.
så
att
Kronan
och
Riddarskapet
näppeligen
tillhopa
har
här
i
Riket
tredjeparten
emot
det
Präster
och
Munkar
/
Kyrkor
och
Kloster
har
.

Väl
bekänner
h
.
N
.
att
han
låter
predika
rena
Guds
ord
och
Evangelium
/
det
vår
Herre
själv
befallt
har
/
och
har
bjudit
samma
predikare
till
svars
/
det
Kyrkans
prelater
icke
har
velat
här
till
dags
undergått
/
utan
säga
att
de
vilja
bli
vid
deras
gamla
sedvänjor
/
evad
hon
är
rätt
eller
orätt
/
emedan
ligga
lekmän
under
och
försvagas
dagliga
dags
mer
och
mer
.

Förs
och
h
.
N
uppå
att
han
vill
inga
Präster
skola
vara
i
landet
/
det
så
uppenbarligen
ljuger
på
h
.
N
.
att
de
som
sådant
utföra
må
sig
skämma
både
för
Gud
och
människor
.

h
.
N
.
akter
dö
en
Kristlig
Man
och
vet
väl
att
vi
icke
kunna
vara
utan
lärare
och
Kyrkopräster
de
oss
skulle
lära
Guds
ord
/
vilka
Lärare
eller
Kyrkopräster
h
.
N
.
vill
styrka
i
all
den
del
de
är
rätta
till
/
så
framt
de
göra
deras
ämbete
fullt
/
det
vet
h
.
N
.
väl
att
man
dem
icke
kan
vara
förutan
efter
skrifterna
/
men
om
de
andra
/
som
det
ämbete
icke
bruka
eller
icke
är
de
meneman
till
tjänst
/
vill
h
.
N
.
veta
ert
goda
råd
/
hur
man
skall
hålla
med
dem
/
efter
i
skrifterna
icke
finns
att
man
dem
behöver
.

Har
och
vår
nådige
Herre
överlagt
sina
uppbörd
och
sina
utgift
och
finns
uppbörden
i
vissa
näppliga
ränta
till
XXIIII.m
.
mark
/
och
utgiften
väl
till
LX.m
.
mark
/
som
h
.
N
.
låter
Er
väl
själva
se
hans
räkenskap
/
och
där
är
med
järnet
inräknad
för
L
.
Lesther
Item
:

Om
det
rop
som
de
har
om
Grijpsholm
.
etc.
kunna
de
icke
annat
säga
/
än
h
.
N
.
är
där
näste
arvingen
till
/
vill
där
någon
om
ropa
vilja
de
var
i
sin
stad
göra
H.N:des
ursäkt
/
och
säga
dem
att
h
.
N
.
är
överbodig
där
om
svarar
varje
och
en
till
rätta
/
och
synes
dem
rätt
vara
att
andra
som
där
till
givit
hade
/
gå
till
rätta
arvingar
igen
/
pantat
och
köpt
löses
till
rätta
börd
.

Och
till
Kronans
upprättelse
efter
hon
försvagat
är
som
h
.
N
.
klagar
/
synes
dem
detta
för
ett
råd
/
att
för
det
rop
skull
som
uppkommit
är
på
Biskoparna
/
att
de
förmäktiga
är
/
så
att
de
Herrar
och
Furstar
i
fordom
har
drivit
av
Riket
/
som
h
.
N
.
klagar
/
må
så
skickas
att
de
skola
över
ens
varda
med
h
.
N
.
hur
mäktiga
H
N
vill
dem
ha
Ridandes
/
vad
sedan
över
är
i
deras
räntor
/
det
skola
de
giva
h
.
N
.
uti
ett
stycke
penningar
efter
som
de
kunna
med
h
.
N
.
över
ens
varda
/
och
h
.
N
.
håller
där
själv
folk
utav
/
och
anammar
till
sig
deras
Slott
besynnerliga
till
dess
Kronans
Slott
/
som
nu
förfallen
är
kunna
igen
uppbyggd
varda
/
och
så
blir
all
for:da
fara
tillbaka
.

Hoppas
Riddarskapet
i
så
måtta
vara
botade
de
drister
som
h
.
N
.
förtält
har
i
sina
framsättningar
/
och
bedja
h
.
N
.
för
Guds
skull
/
att
han
dem
icke
än
nu
utöver
giver
/
utan
blir
vid
Riket
styre
och
råd
som
här
efter
som
här
till
dags
/
de
vilja
vara
h
.
Nådes
Tro
män
/
i
döden
där
skall
h
.
N
.
förlåta
sig
uppå

Efter
Clerkerijd
är
och
en
stor
sack
där
till
ju
en
part
av
dem
/
må
allvarliga
sägas
Kyrkans
prelater
till
att
de
sådana
avstilla
med
sina
Klerker
/
eller
dem
skall
därom
tilltalas
som
deras
Klerker
bruka
/
och
att
sådana
skall
varda
strafat
vilja
alla
Köpstädesmän
tillhjälpa
med
liv
och
makt
;
Det
samme
säljs
och
fogdar
/
Borgmästare
och
Råd
i
städerna
allt
de
sådana
stämplare
straffa
där
de
dem
förnimma
/
eller
svarar
de
där
till
.
etc.
Item
:

Om
denne
nye
tro
eller
lärdom
som
sägs
vara
uppkommen
nyligen
här
i
Riket
/
är
väl
sant
att
mycket
fåfängt
ryktas
därom
/
som
munkar
och
präster
har
oss
föregivit
/
dock
efter
det
övergår
vårt
föga
förstånd
skjuter
vi
det
in
till
de
goda
män
som
Höglärda
och
i
skrifterna
väl
förfarna
är
/
vilka
som
ytterligare
där
om
rannsaka
kunde
/
som
är
Bispar
/
Prelater
.
etc.
att
de
ville
granneliga
överväga
vad
rätt
eller
orätt
var
/
begärandes
för
den
skuld
högeliga
av
vår
K
.
N
.
Herre
/
att
H
,
N
.
ville
låta
komma
dem
tillhopa
som
denne
sack
mest
anrör
i
vår
närvaro
/
så
att
vi
måtte
bli
rätteligen
undervisade
i
det
som
rätt
och
kristligt
vore
.

Den
första
för
den
ostadighet
skull
som
plägar
vara
i
Riket
/
den
h
.
N
.
och
befunnet
hade
i
sin
tid
med
många
stämplingar
och
uppstöter
/
som
emot
H
N
.
skedda
vore
/
som
var
av
Herr
Pedher
Canceller
och
hans
parti
och
nu
med
den
förrädare
i
Dalarne
/
som
sig
kallar
h
.
Stens
Son
/
av
vilka
vill
efterfölja
att
om
några
ville
sig
företaga
något
obestånd
i
Riket
/
behöver
han
ej
annat
göra
än
giva
sig
tid
upp
/
och
då
har
man
strax
uppenbarlig
orligh
och
obestånd
/
för
vad
sack
dem
själva
täckes
föregiva
sann
eller
osann
/
och
bli
slika
skalkar
och
stämplare
där
och
annorstädes
i
landet
så
betrodda
att
de
må
dristeliga
och
ostraffad
säga
på
h
.
N
.
och
på
vem
dem
!
täcks
allt
det
dem
lyster
och
har
för
den
skuld
alla
de
som
förräderi
har
i
sinnet
eller
de
som
åstunda
till
Riket
inländska
eller
utländska
god
råd
där
med
fullfölja
deras
uppsåt
och
mening
:

Och
hade
h
.
N
.
samma
predikare
till
städes
och
bjöd
dem
till
svars
om
där
några
hade
varit
av
Clerkerijd
som
dem
hade
velat
tilltala
och
vinna
dem
till
några
oredliga
stycken
i
deras
lärdom
/
var
så
skedde
ville
h
.
N
.
då
straffa
dem
/
som
tillbörligt
vore
/
var
och
icke
/
begärde
då
h
.
N
.
att
vi
råd
skulle
finna
emot
för:ne
rop
/
såsom
på
h
.
N
.
orätteliga
påfördes
.

Till
att
bota
den
första
bristen
/
lovade
vi
h
.
N
.
som
vi
och
med
detta
vårt
öppna
brev
lovar
vid
vår
ära
och
redlighet
/
var
i
sin
stad
/
vilja
hjälpa
till
att
straffa
de
slika
rop
/
rykte
/
och
obestånd
åstad
komma
emot
h
.
N
.
evar
det
helst
ske
kan
i
Dalarna
eller
annorstädes
/
och
så
bevisa
oss
med
h
.
N
.
att
i
de
måtten
näst
Guds
hjälp
ingen
fara
skall
vara
till
någon
förvandling
i
Riksens
regemente
antingen
för
utländska
eller
inländska
.

Vi
Gostaff
etc.
hälsar
Er
tack
vi
Er
alla
kärliga
för
Er
godvillighet
/
hulskap
/
troskap
och
lynne
som
I
oss
i
alla
måtte
troliga
bevisat
har
;
och
änkannerliga
nu
med
denne
utgjorda
Giärd
och
hjälp
till
Riksens
gälds
betalning
/
därför
vi
gärna
vilja
veta
ert
bästa
.

För
Hor
/
Lönskeläije
,
Jungfrukränkning
/
bötas
Konungen
och
icke
Biskopen
.

Där
Präster
eller
Lekman
stå
var
annan
/
vare
icke
den
ena
mer
i
Ban
än
den
andra
/
efter
Gud
har
så
väl
förbjudit
den
ena
slå
som
den
andra
/
utan
bötar
var
för
sin
Sak
efter
Landslagen
.

Vi
befaller
och
Lands
och
Fjärdingsmän
att
de
är
dem
med
Skjutshästar
och
all
annan
nödtorftig
fri
fordenskap
beforderliga
så
länge
denne
rannsakning
uppå
står
där
var
och
en
i
sin
stad
som
för
vår
skull
ville
och
skola
göra
och
Låta
veta
sig
hörsamligen
efter
rätta
,
av
Gripzholm
den
6
februari
år
1622
.

Vorde
Morthen
och
Olof
förenade
och
Lades
40
daler
i
vi
de
den
sig
på
den
andre
först
förbryter
.

Olof
,
Arfwedz
dräng
i
Vmberga
hade
gjort
mökränkning
med
Jngel
barn
född
i
Danmora
Socken
vart
sack
40
mr
.
lyftesmän
Per
Joensson
i
Anebo
.
h
.
Valborg
drängens
Styvmoder
drängen
tjänar
nu
på
Öreby
och
skall
ha
för
sin
tjänst
av
Sonen
10
daler
.

Sockenstugan
Närvarandes
Kronans
befallnings
Man
,
där
samme
städes
Ärlig
välaktad
och
förståndig
Oluf
Jönnssonn
dessa
Ärligen
Edsvor
,
Danne
mäns
satt
i
Nämnden
,
Hans
Larssonn
i
öster
Ekeby
Matz
Anderssonn
ij
Kålboo
do
:

Lars
Andersonn
i
w
Ekeby
Tomas
Matzonn
i
Grythby
Oluf
Andersonn
i
Bökreby
Lars
Andersson
i
Brunby
Samma
Dag
Kom
för
rätten
hans
Abrahamsonn
i
Skarp
Ekey
och
På
av
beredde
mode
och
god
vilja
såsom
och
med
sin
hustrus
broder
Ja
och
Samtycke
sålde
och
upplät
hustru
Anna
i
jerssmyra
all
den
arv
del
Dem
till
fallit
var
uti
be:te
Jerssmyra
och
där
förre
uppbör
nu
strax
reda
Penningar
25
daler
och
i
Vängåvor
en
sked
om
tre
Lod
,
Där
om
de
nu
vorde
vänligen
och
väl
förlikta
och
gjorde
var
andra
hade
sträckning
in
för
sittande
rätten
Så
alldenstund
detta
köp
Lagligen
gjort
var
såsom
och
Lagbudet
och
Lagståndet
,
som
Lag
före
Dömde
och
ingen
nu
var
som
här
å
talade
eller
tala
ville
,
där
för
Dömde
iag
samt
Nämnden
Detta
köp
Stadigt
och
fast
att
Stånda
och
aldrig
återigen
här
å
tala
vid
vars
och
3
mr
förhärdsdöm
S
D
Var
Pedirr
Andersonn
i
trosberg
Stämd
av
Nämndeman
att
Svar
Befallningsmannen
kom
in
:
tillstädes
vart
därför
saker
till
3
mr
till
vidare
rannsakning
.

Vart
allmogen
förmanad
att
när
de
få
bud
skola
de
komma
vid
bot
[
Lars
Erichsson
i
Abyggeby
blev
tilltalad
på
Hans
Larssons
en
borgares
i
Gäfle
vägnar
om
i
t:na
korn
då
sade
han
att
h
.
Olof
i
Thensta
hade
tagit
samma
korn
t:na
för
det
Hans
var
honom
skyldig
2
t:nor
krampsill
,
vart
sagt
att
Lasse
skulle
betala
Hans
och
Lasse
gå
till
Prästen
.
]
5
Olof
Persson
i
Hwseby
hade
löpt
efter
sin
Stiufsson
Erich
Olofsson
i
Hökeby
in
till
hans
gård
och
slagit
på
hans
port
med
en
stör
,
som
han
icke
kom
in
ville
han
kliva
över
balken
in
till
honom
,
och
då
ingen
mera
skada
gjorde
vart
sak
för
hemgången
40
mr
.

(
1631
)
Den
31
Januari
stog
Lagting
uti
Befallningsmannens
Ärlig
och
välaktat
Hans
Larssons
närvaro
dessa
Edsvurna
satt
i
Nämnden
.

Noch
frikallades
h
.
Brijta
i
Westerijcke
för
h
.
Margretas
i
Torkilsboo
i
Wendels
Socken
ogrundade
tillmäle
som
dock
där
om
ingen
skäl
eller
liknelser
finnas
kunde
,
och
Sattes
därhos
vite
att
hon
henne
här
Utinnan
ytterligare
vräker
skall
vara
Sacher
till
Penningar
-
40
mr
.

Item
tillsades
efter
hennes
M:tz
vår
allranådigaste
Drottnings
brev
,
att
alla
skola
sig
vargnät
förskaffa
.

Noch
vittnade
och
bekände
Nämndemännen
att
Peder
Larsson
i
Bålemyre
,
hade
nästförlidna
höst
som
var
S
Mathias
afton
,
igenom
häftig
vådeld
,
bortmist
först
både
man
och
Ladugård
,
att
icke
en
husknut
är
kvarbliven
:

Noch
vittnade
Nämnden
att
de
två
öres
Land
Kronojord
i
Läby
Uti
Biorklinge
Socken
,
sm
nu
där
sammastädes
hävdar
och
brukar
,
kunde
inte
:
göra
skäl
för
'
/
»
Mantal
,
och
fördenskull
där
th
:
icke
kunde
Uti
*
/
4
hemman
förmedlas
,
blir
det
och
alldeles
öde
.

Alltså
visste
icke
härads
Nämnd
hans
Liv
i
Någon
måtto
att
befria
,
och
fördenskull
Såsom
han
människo
blod
Utgutit
har
:

Vart
sagt
att
Syn
skulle
dit
och
där
om
granneligen
rannsaka
med
det
förste
.

Köpslog
och
Lars
Joensson
med
sin
Syster
dotter
fönne
h
.
Brita
om
hennes
del
i
Jord
och
hus
i
Grimsarebo
och
vorde
således
för
enade
att
Lasse
skulle
giva
henne
till
den
Silverkosa
hon
bekommit
hade
Spannmål
2
t:nor
,
där
på
de
gjorde
var
andra
handsträckning
.
fönne
Jord
uppbjöds
förste
sin
.

Morthen
Persson
i
Österekeby
Hans
Humbla
i
Äkra
.
domare
Lars
Andersson
i
Westerekeby
Lars
Andersson
i
Brunby
Matz
Andersson
i
Kårbo
Thomas
Matsson
i
Grytteby
Erich
Staphansson
i
Tolsmyra
(
Arfwedh
Persson
i
Vmberga
)
(
Erich
Håkansson
i
Grytteby
)
Nils
Persson
i
Äkra
lät
tredje
sin
uppbjuda
det
hemman
han
besitter
och
köpt
hade
av
sina
Syskon
som
är
Lars
och
Per
Perssöner
.
h
.
Anna
i
Karby
h
.
Elin
i
Skarpekeby
(
och
dem
betalt
)
.

Befallningsmannens
välbetrodd
Anders
Hööck
besvärade
sig
att
ha
låtit
uppbära
någon
humbla
och
fläsk
med
ett
Betzman
som
ringare
är
på
vart
få
till
2
mr
som
Proberat
var
här
för
rätten
och
fälldes
efter
det
rätta
betzmannet
,
och
var
kommen
till
korta
på
humblan
i
få
16
mr
vart
sagt
att
den
som
hade
levererat
med
den
ringa
vikten
skulle
betala
det
som
felar
(
h
.
Jngri
i
Alderbecken
besvärade
sig
att
det
fordras
av
henne
Qwarntuls
Mantals
Penningar
för
den
dräng
hon
hade
stått
sig
och
sedan
låtit
Lägga
sig
till
knekt
av
Lars
Morthensson
i
Ekeby
,
vart
sagt
att
Lasse
där
han
är
skall
betala
för
honom
de
6
mr
som
skall
Låta
malå
för
honom
)
Wendel
och
Börklinge
Socken
:

Då
ropade
Erich
och
sade
,
kör
intet
hit
,
Jag
fruktar
träd
faller
,
övergav
så
Erich
att
hugga
då
körde
Andes
till
sin
stock
,
när
han
hade
vänt
kälkarna
till
,
och
skulle
Lassa
uppå
föll
träd
om
kull
och
in
på
Andes
att
han
blev
där
död
Liggande
.
(
Som
och
S
.
Anders
Larssons
Son
som
med
var
i
skogen
berättade
,
som
och
Olof
och
Thomas
i
Husby
vittnade
som
och
där
vore
)
Vart
Erich
sack
efter
det
9
Kap.
i
dråp
:

Vart
sagt
att
Per
skulle
giva
14
daler
igen
,
då
vorde
de
så
överens
att
Erich
skulle
ha
ett
Äng
som
Räntar
4
lass
hö
om
året
till
dess
han
bekommer
sina
Pengar
igen
,
dock
skulle
det
vara
gott
slags
hö
.
(
h
.
Brita
And
ers
Anderssons
i
Tolbon
i
Börklinge
Socken
kärade
till
Jahan
Orm
i
Klarengie
om
4
daler
12
öre
kopp:mynt
där
på
hon
hade
uppburit
en
halvspann
Råg
för
6
mr
Resterar
henne
2
daler
28
öre
,
lovade
betala
innan
14
dagar
vidare
bot
.

Då
kom
för
rätten
den
Ädel
och
välboren
Frues
Fru
Christinas
Sigri
Bielkes
till
Öreby
Predikant
välLärd
h
.
Abraham
och
på
Hennes
N:s
vägnar
böd
efter
fönne
hemman
medan
h
.
N:d
tilkommer
årlig
skatten
(
och
utlagorna
)
efter
bytes
brevet
och
Adliga
Privilegier
vara
tet
Närmast
,
sköts
upp
att
vidare
(
förskaffa
)
hos
höge
över
heten
(
brev
därpå
,
medan
Lars
Andersson
hade
det
köpt
,
sedan
det
var
h
.
N:d
tillbudet
,
och
h
.
N:d
icke
hade
givit
där
Guds
Penning
på
)
.

Oloff
Matzsson
i
Skarpekieby
lät
annat
sin
uppbjuda
det
hemman
han
besitter
och
köpt
har
av
sina
systrar
och
syster
barn
[
Befallningsmannen
befallde
och
tillsade
allmogen
som
pläga
bygga
vägen
här
ifrån
Socknen
,
och
till
Tegelsmora
att
de
den
med
det
första
förfärdiga
att
han
blir
laggill
och
god
vid
straff
.
]
3
Hederligh
och
välLärd
h
.
Anders
Prost
och
Kyrkoherde
i
Wendel
Socken
lät
förste
sin
uppbjuda
sitt
och
sin
S
.
Broders
Staphan
Erssons
(
bars
)
hemman
i
Berghby
,
som
wälbe:te
Herr
Andersses
inlagda
skrift
i
Rätten
vidare
förmäler
Marten
Persson
i
osterekieby
dorn
Matz
Hansson
i
Grytby
Hans
Humbla
i
Äkra
Lass
Persson
i
läby
Lass
Matzsson
i
Osterekieby
Lass
Andersson
i
Westerekieby
Matz
Olofsson
i
Kaslinge
Arfue
Persson
i
Vmberga
Erich
Staphansson
i
Torsmyra
Öffersten
Ädel
och
välbördig
Mauritz
Magdual
till
broby
berättade
att
hans
Syster
hade
insänt
en
Tysk
Fänrik
att
utfordra
någon
gall
,
som
de
har
att
fordra
efter
sin
S
.
Moder
,
så
emedan
deras
S
.
Moder
är
än
obegraven
och
efter
hennes
begravning
skifta
arvet
.

Ävenledes
hade
gruvfogden
Johan
Upström
instämt
torparen
Olof
Halfwarsson
i
Stenstugan
för
en
skuldfordran
av
43
daler
kopparmynt
,
men
gav
till
känna
,
att
de
för
denna
gången
sålunda
överens
kommit
,
att
svaranden
skall
sig
hos
käranden
infinna
och
därom
göra
behörig
räkning
;
Varför
ock
rätten
lämnade
det
där
vid
till
vidare
.
/
Gruvfogden
välbetrodde
Johan
Uppström
hade
också
instämt
bonden
Anders
Andersson
i
Fåneby
för
en
skuld
fordran
av
45
daler
kopparmynt
samt
och
Anders
Pehrssons
arvingar
i
Brunby
för
16
daler
16
.
/
.
kopparmynt
,
vilka
summor
han
påstått
att
få
befallde
jämte
expenser
,
men
gav
nu
för
rätten
till
känna
,
vad
den
förra
eller
Anders
Andersson
angår
,
det
de
med
var
annan
därom
sålunda
kommit
överens
och
till
förliknings
,
att
Anders
Andersson
skall
i
ett
för
allt
till
honom
betala
24
daler
kopparmynt
;
och
vad
Anders
Pehrssons
arvingar
i
Brundby
beträffar
,
så
emedan
mågen
Erich
Ohlsson
berättade
,
att
herrskapet
tagit
av
dem
allt
det
de
hade
efter
bemälde
Anders
Pehrsson
för
skuld
,
vilket
ock
nämnden
med
flera
närvarande
intygade
;
Ty
gav
Upström
denna
sin
fordran
efter
,
var
vid
fördenskull
rätten
lät
bero
och
förbli
.
/
Befallningsmän
herr
Philip
Befvert
på
Kiettslinge
hade
väl
instämt
tolvmannen
Erich
Ersson
i
Råmstarbo
för
den
ohägn
och
skada
en
hans
häst
skall
gjort
honom
på
Kietzlinge
tillhörige
äng
i
Karboda
,
varför
han
påstått
laga
plikt
,
skadans
ersättning
jämte
expenser
,
men
gav
för
rätten
tillkänna
,
att
Befvert
sådant
eftergivit
och
lämnat
,
emot
det
att
Erich
Ersson
skall
hjälpa
honom
något
,
när
han
litar
honom
till
;
Ty
lämnade
rätten
det
där
vid
.

Jan
Ersson
tillspordes
alltså
,
varifrån
han
fått
anledning
till
att
således
stämma
denna
sin
hustru
?

Karin
Erichsdotter
,
efter
stämning
tillstädes
,
tillstod
,
att
hon
så
sagt
och
att
det
är
sant
,
det
hon
,
om
så
skulle
behövas
,
med
vittnen
skall
kunna
bevisa
,
men
om
de
bedrev
någon
otukt
med
var
annan
,
sade
hon
sig
intet
veta
eller
kunna
säga
.

Hoffman
,
att
emedan
denna
gärds
gård
intet
hör
StorEnen
utan
Norrby
till
,
så
vill
man
vidare
svara
här
till
,
när
man
å
Norrby
sida
blir
därom
lagligen
stämd
och
tiltalad
.

Anno
1736
den
32
och
4
maj
hölls
ordinarie
laga
sommarting
med
allmogen
och
menige
man
av
Wändels
socken
och
tingslag
,
närvarande
Kronans
länsman
välaktad
Gabriel
Wretberg
och
tingslaget
vanliga
och
nedanskrivna
nämnd
,
nämligen
:

Och
jag
,
Erich
Boije
,
där
emot
uppdrager
till
herr
löjtnant
Pehr
Pehr
Leufstedt
mitt
halva
hemman
,
Kullbohl
benämnt
,
/
med
allt
vad
samma
hemman
tillkommer
,
såsom
jord
,
hus
,
etc
,
intet
undantagande
,
samt
och
även
lämnat
och
betalat
och
betalat
till
herr
löjtnant
Leufstedt
,
såsom
en
mellangift
på
detta
oss
emellan
skedde
byte
,
tvåtusende
daler
kopparmynt
,
vilka
2000
daler
,
den
första
penningen
med
den
sista
,
såsom
jag
,
Pehr
Leufstedt
,
redan
av
kyrkoherden
handfånget
,
ty
skall
ock
detta
byte
fast
stånda
och
icke
något
klander
och
åtal
på
någondera
sidan
av
oss
,
under
vad
pretext
det
vara
kunde
,
vidare
här
på
göras
,
kommande
vi
nästkommande
Tomassmässo
våra
bönder
på
samma
våra
hemman
att
lagligen
uppsäga
och
,
sedan
de
sin
laga
f
ardag
njutit
,
till
varandra
samma
hemman
,
som
ovanförmält
är
,
att
avträda
.

Nils
Pärsson
kom
intet
tillstädes
utan
berättades
av
länsmannen
vara
utur
socknen
bortgången
,
utan
att
han
vet
,
varest
han
nu
är
tillfinnandes
.

Responsum
,
att
klockan
kunde
vara
10
om
aftonen
.

Vad
utsädet
anbelangar
,
så
tillstod
Brundin
,
att
han
fått
3
tunnor
om
året
av
råg
,
korn
,
havre
och
blandsäd
till
att
så
ut
på
Ohsengii
halvdel
samt
att
det
så
gått
till
,
att
han
undertiden
har
måst
lägga
mera
därtill
.

Ekeroth
tillstod
detta
så
,
att
han
gick
till
Håfgårdzberg
emellan
predikningarna
och
köpte
för
3
.
/
.
brännvin
,
till
förekommande
att
sjukdomen
,
varav
han
under
ottesångspredikan
skall
haft
starka
känningar
,
intet
måtte
taga
överhanden
hos
honom
.

Quasstio
,
hur
länge
han
varit
under
krigstjänsten
?

Uti
den
av
Bängdt
Bängdtsson
i
SkarpEkeby
emot
Anders
Ersson
i
Smedby
instämde
sak
om
en
skuld
fordran
av
48
daler
kopparmynt
och
1
/
2
tunna
råg
,
dem
han
påstått
att
få
jämte
intresse
och
expenser
befallde
,
angav
de
sig
sålunda
vara
förlikta
och
överens
komna
,
att
Bängdt
Bengtsson
fått
4
plåtar
av
svaranden
och
att
han
inom
2
år
skall
få
två
plåtar
till
samt
få
,
för
det
han
väntat
och
för
sitt
besvär
,
slå
en
äng
till
3
lass
i
två
år
Mårten
Mattsson
i
Allerbäcke
hade
väl
instämt
Anders
Pehrsson
i
Tråtzberg
angående
en
bössa
,
som
Anders
Ersson
/
skall
av
Mårten
Mattsson
lånat
,
och
fördenskull
påstått
att
få
igen
jämte
expenser
,
men
gav
nu
tillkänna
sig
sålunda
vara
därom
förlikta
och
överens
komna
,
att
käranden
lämnat
svaranden
tid
till
nästkommande
kyndermässa
att
skaffa
bössan
igen
,
vilken
skall
blivit
för
honom
bort
stulen
,
och
där
hon
då
intet
kan
fås
igen
,
skall
han
betala
henne
med
tolv
daler
kopparmynt
;
fördenskull
lät
rätten
det
därvid
bero
och
förbli
.

Men
Svinhufwud
sade
sig
ingen
stämning
härom
ha
fått
,
som
han
icke
heller
för
den
,
utan
för
annan
orsak
kommit
hit
till
tinget
.

Och
som
Råkne
,
sedan
han
av
Hagels
bok
blivit
underrättad
,
varuti
skulden
består
,
den
intet
gitte
disputera
,
/
och
han
så
väl
som
Hagels
fullmäktig
,
dess
son
gruvfogden
välbetrodde
Carl
Hagel
,
var
nöjda
där
med
,
att
denna
Råknes
skuld
skall
,
efter
befallningsmannen
välbetrodde
Philip
Befwerts
nu
här
in
för
protokollet
givna
försäkran
,
bli
för
Råkne
betalat
vid
Leufsta
bruk
;
Så
lät
ock
rätten
det
där
vid
bero
,
och
prövades
för
övrigt
skäligt
,
det
bör
Råkne
dessutom
uti
expenser
till
inspektorn
Hagel
erlägga
sina
6
daler
kopparmynt
.

Matts
Andersson
i
Åhl
,
som
av
inspektorn
herr
Erich
Hagel
var
instämd
om
24
daler
24
.
/
-
kopparmynts
skuld
,
förnams
vara
sjuk
och
hade
således
laga
förfall
,
varför
som
Hagells
fullmäktig
förbehöll
sig
att
få
vid
nästa
ting
tala
honom
härom
till
,
så
stannade
det
där
vid
för
denna
gången
.

Däremot
sökte
Erich
Ersson
att
försvara
sig
med
en
den
7
angusti
1682
emellan
Frebro
och
Fastebo
i
Tiärp
av
lagläsaren
Matthias
Erling
och
Tiärpz
härads
nämnd
in
loco
förrättad
rågång
syn
,
varav
fanns
,
att
Barsmosse
och
Kohlswedzrören
blivit
erkända
för
rätt
skillnad
på
södra
sidan
emellan
Frebro
och
Fastebo
,
vilket
ock
fanns
vara
vid
tinget
år
1683
den
11
oktober
uppläst
och
konfirmerat
.

Johan
Andersson
tillstod
,
att
han
huggit
7
stycken
klabbar
på
allmäningen
,
allenast
sex
å
7
alnar
långa
,
men
ville
ursäkta
sig
där
med
,
att
han
såsom
nyss
kommen
till
Botarbo
intet
visste
,
huruvida
Botarbo
ägor
sträcka
sig
utom
deras
odal
hank
och
stör
.

Länsmannen
beropade
sig
alltså
på
sina
instämda
vittnen
Anders
Ersson
i
Giärsmyra
och
klockaren
Jan
Ersson
,
vilka
ojävade
avlade
vittneseden
och
berättade
var
för
sig
,
först
Anders
Ersson
,
att
han
såg
,
det
Anders
Olssön
då
var
drucken
;
men
Jan
Ersson
,
att
han
det
intet
såg
utan
kunde
allenast
så
tycka
,
eftersom
han
sätt
och
kved
vid
bordet
,
varför
de
andra
hade
honom
ut
,
på
det
han
intet
måtte
förarga
herr
kyrkoherden
;
I
anseende
var
till
,
och
emedan
allenast
det
ena
vittnet
sett
honom
,
Anders
Olssön
,
den
gången
vara
drucken
,
men
det
andra
intet
,
han
från
länsmannens
tilltal
härom
befriad
varder
,
i
följe
av
Kungl.
Maij:ts
nådigaste
plakat
om
svalg
och
dryckenskap
av
år
1733
och
dess
2

Land
ägaren
välbetrodde
Anders
öhrling
hade
också
låtit
inkalla
följande
för
försummat
drevskall
till
björnars
uppletande
nästlidna
den
3
,
4
och
5
januari
,
nämligen
Åkra
gamle
Michel
Ersson
,
Huseby
Michel
Ersson
,
Falsboda
Matts
Mattsson
,
Bärgby
sergeanten
Elgklo
,
ibidem
Pär
Pärsson
,
Kietzlinge
befallningsmannen
Philip
Befwert
,
Ängen
Erich
Ersson
,
Grytby
Anders
Jacobsson
,
Kläringe
Olof
Jansson
,
Gulboda
Olof
Ersson
,
Slubolet
Olof
Ersson
och
Råssla
Jan
Pärsson
;
men
som
det
befanns
,
att
de
alla
hade
laga
förfall
,
i
det
de
dels
vore
borta
,
när
skallet
blev
pålyst
,
dels
sjuka
och
ensamma
karlar
,
när
det
stod
,
dels
torpare
under
säterierna
Öhrby
och
Kietzlinge
,
från
vilka
alla
deras
övriga
torpare
,
när
Olof
Jansson
i
Ängen
,
Olof
Ersson
i
Slubolet
och
Jan
Pärsson
i
Råssla
då
vore
sjuka
,
bevistat
detta
skall
;
Ty
blir
de
från
böter
denna
gången
befriade
.

Följande
har
vid
detta
ting
begärt
timmer
och
byggnings
virke
samt
gärdsel
och
stor
efter
vederbörlig
skedde
syner
och
besiktningar
,
nämligen
'
:

Upplästes
landshövdingens
välb:
Hans
Strijks
brev
,
angående
den
skuld
och
rättighet
som
Elin
Kruse
har
att
fordra
på
sin
S
:
förre
mans
Clas
Larsson
lagmanstull
.

I
lika
måtto
har
be:te
Hans
Erichsson
till
fullo
nöje
utbetalt
Måns
Oluffsson
för
en
fjärde
part
och
i
be:te
gård
liggandes
med
30
Rd:r
och
seendes
är
av
deras
gjorda
underskriven
köpeskrift
,
så
att
summan
84
Rd:r
belöper
sig
som
förbe:te
Wästergården
Gränåås
utgiven
är
,
den
siste
med
den
förste
penning
uppburen
och
riktigt
betalat
har
.

Samma
dato
anpresenterade
ärlig
och
beskedlige
danneman
Erik
Olofsson
,
ett
lagbudet
och
ståndet
köpebref
där
med
bevisandes
sig
lagligen
ha
köpt
Jonsgården
av
Erik
Persson
ibidem
;
Och
nu
därför
levererat
allra
först
till
hans
åtskilliga
kreditorer
fyrtio
Rd:r
såsom
och
givet
för
ett
genlagt
pantgods
och
åkerstycke
kallat
Brodswedh
elva
Rd:r
,
blir
alltså
summan
femtio
och
en
Rd:r
,
vilket
köpebrevet
och
med
följande
specifikation
bredare
utvisar
.

Anklagades
ryttaren
Hindrik
Hyldh
vilken
mökränkning
gjort
med
en
jänta
Elin
Eriksdotter
i
Sikås
,
varför
rätten
honom
tillsporde
om
han
detta
gjort
har
,
var
till
han
sig
skyldig
gav
,
men
sade
sig
henne
inte
något
äktenskap
ha
lovat
.

(
2
)
Länsman
Claes
Isaksson
Kiock
angav
i
Rätten
det
Anders
Jönsson
i
Strand
,
har
hyssat
2:ne
förrymde
ryttare
,
nebl:n
fan
junkaren
Per
Jönsson
som
för
några
år
sedan
utan
någon
orsak
rymde
,
undan
welb:n
H
Ryttmästarens
Gerhardt
Gernfeldts
kompani
till
Norge
där
han
allt
härtill
har
tillhållit
,
men
nu
åter
rymt
från
Norrighe
havandes
med
sig
i
följe
en
Norriges
korpral
,
Anders
Skåningh
som
tillika
med
sin
hustru
har
där
ifrån
rymt
och
begivit
sig
utför
åt
Ångermanland
,
och
omsider
nu
epargeras
,
att
dessa
har
stulit
i
Norrige
en
stor
post
penningar
,
och
sedan
rymt
där
ifrån
vilka
har
kommit
till
Ströms
s:n
,
hos
denne
Anderss
Jönsson
i
Strand
och
begärt
hus
om
natten
hos
honom
,
vilket
han
dem
ej
förvägra
kunde
,
utan
skickade
genast
efter
förridaren
under
dragonerna
,
Olof
Jonsson
Klöster
,
i
den
mening
att
förhöra
vad
det
skulle
vara
för
ett
parti
efter
de
reste
så
Fjäll
vägen
,
och
sedan
skulle
han
med
sina
dragoner
dem
fast
taga
,
vilket
Olof
Jonsson
ej
efterkom
;
utan
förblev
hos
dem
och
Förridaren
kände
Fanjunkaren
igen
som
här
från
Jemptelandz
Kompani
förrymd
var
,
men
ingen
tog
honom
fast
,
utan
lät
dagen
efter
fara
dem
sin
väg
.

(
18
)
Dessutom
har
denne
lapplandsman
Lars
Larsson
hyst
och
undan
dolt
en
norriges
lap
,
Thomas
Persson
som
har
rymt
från
Norrighe
och
icke
uppenbarat
för
befallningsman
då
han
kom
till
honom
i
fjället
för
än
de
andra
angav
honom
.

(
21
)
Kyrkoherden
i
Hammerdahl
well:de
H:r
Erik
Hedsander
,
äskar
och
begär
syn
nästkommande
sommar
,
emellan
sig
och
sina
grannar
Måns
Eriksson
i
Mo
,
och
Lars
Persson
i
Bye
angående
kyrkomyran
;
Såsom
och
ett
prov
och
rann
sakning
på
hans
skog
och
slott
,
och
emedan
som
en
av
konsistoriets
wäg:r
bör
tillstädes
vara
,
ty
bör
kyrkoherden
angiva
sådant
hos
h:s
vördighet
Prosten
.

Olof
Eriksson
i
Ede
Anders
Sjulson
i
Fyrås
Per
Danielsson
i
Grelsgård
Nils
Andersson
i
Tullingsås
Christen
Persson
i
Viken
Olof
Andersson
i
Solberg
Jöran
Andersson
i
Öhn
Erik
Samuelsson
i
Håxås
Per
Broddesson
i
Öhn
Nils
Andersson
i
Ede
Per
Eriksson
i
Sikås
Olof
Thorsson
i
Hallen

Måns
Eriksson
i
Mo
låter
uppbjuda
sin
gård
andra
gången
,
nästa
frände
tillåter
lösen
.

B
.
och
där
på
befallningsmannens
wälb:de
Daniel
Bertilssons
kvittens
på
det
ena
1660
års
resterande
ödes
utlagor
,
som
dokumentet
lit
C
.
de
dato
Mo
28
November
1666
förmäler
var
av
sedan
följer
Anders
gården
vara
efter
H:s
Excell:tz
Guvernörens
restitution
till
odel
kommen
,
ödes
utlagorna
betalade
blev
.

Kap.
Ärvde
ballken
har
sig
regulerat
och
sökt
sin
arvs
pretension
innan
\
natt
/
jämn
långa
,
var
ifrån
denne
Rätten
ej
kan
gå
,
utan
stadig
hålla
sig
där
vid
;
berörde
odelsmän
det
samma
icke
allenast
försuttit
,
utan
för
14
.
år
sedan
från
Jemptelandh
sig
begav
och
sitt
odels
hemman
övergav
,
var
igenom
det
är
blivet
öde
och
kommit
till
stort
van
bruk
,
Kronan
och
dess
boende
till
ingen
ringa
kostnad
,
allt
där
före
resten
6½
Rd:r
Kronan
tillkommer
som
bemält
är
,
belöper
Summan
27
.

LL
och
söker
sin
man
,
det
bäst
de
gitta
,
Jemptskogswägen
allenast
angående
.

Men
intet
nedersätta
sig
någorstädes
till
annans
förfång
eller
skada
,
som
dels
här
till
skett
är
.

Sammaledes
Olof
Larsson
i
Gåxsjö
skall
och
komparera
på
nästa
ting
,
och
svara
för
det
han
har
varit
borta
på
andra
storböndagen
.

Jon
Sjulsson
i
Vallen
och
Ström
socken
,
som
lagligen
stämd
är
att
svara
till
Olof
Olofssons
pretension
på
en
ök
,
sakfälldes
efter
33
kap.
tingm.b
.
för
stämnings
försittande
3
mk:r
.

Länsman
Christian
Andersson
angiver
det
Lars
Nilsson
i
Nääs
,
har
lägrat
pigan
Gunborg
Jonsdotter
i
Öhn
,
vilket
Lars
tillstår
;
men
Gunbor
för
sitt
sjuklige
barn
och
detta
stora
oföre
ifrån
Ström
socken
,
ej
tillstädes
är
,
ty
uppsköts
detta
till
nästa
laga
ting
,
efter
tolvman
Per
Broddesson
berättar
,
det
Gunbor
har
för
sig
bekänt
att
Lars
har
lovat
henne
äktenskap
.

Emedan
som
Olof
Andersson
i
Solberg
för
rätten
bekänner
och
tillstår
,
ha
uti
3
års
tid
uppgrävt
lönn
gravar
på
kronägorna
som
länsmans
hemmanet
Ede
tilhör
,
och
där
fångat
en
liten
älg
som
han
själv
bekänner
.

Kronans
länsman
Christian
Andersson
angav
i
rätten
ha
förnummit
av
Wellam
Persson
i
Fyrås
förliden
midsommars
dag
1674
,
att
Jöns
Jonsson
och
Jon
Hemmingsson
i
Fyråås
har
uti
förbjuden
tid
afton
för
full
?
)
midsommars
dagen
fört
hem
ur
skogen
en
full
vuxen
älg
,
och
att
de
fjärde
dag
pingst
har
gått
till
skogs
med
bössa
och
2
.
hundar
haft
med
sig
,
förmenar
att
djuret
då
har
blivit
skjutet
,
efter
det
var
allenast
14
dagar
emellan
de
det
hemförde
.

När
de
kom
dit
,
blev
de
intet
något
djur
varse
,
allenast
de
såg
spår
eller
fjät
efter
älgen
,
sedan
föregiva
de
ha
gått
tillbaka
,
då
de
,
under
vägen
mötte
Wellam
Persson
i
Fyhråås
.

Anders
Mårtensson
i
Öhn
,
avlade
sin
nämndemans
ed
.

Och
ehuruväl
på
åtskilliga
Tider
/
och
mest
uppå
alla
Riksdagar
/
vid
pass
50
à
60
År
tillbaka
/
är
vordet
omtalat
och
påmint
/
att
Kyrkobalken
/
och
den
i
trycket
för
detta
utgångna
KyrkoOrdningen
/
skulle
överses
och
förbättras
/
var
till
och
så
åtskilliga
utkast
/
Tid
efter
annan
är
gjorda
;
så
har
likväl
Överhetens
goda
uppsåt
/
och
Undersåtarnas
billiga
åstundan
/
allt
här
tills
stannat
uti
en
ofullkomlighet
/
för
åtskilliga
hinders
skull
/
som
alltid
har
legat
ett
så
viktigt
Verks
fullbordan
i
vägen
.

De
Kristliga
Ceremonier
,
som
här
till
uti
våra
Församlingar
har
varit
i
bruk
/
och
ännu
brukas
/
oansett
de
är
i
sig
själva
villkorliga
/
och
intet
göra
till
Saligheten
/
skola
de
likväl
/
såsom
till
en
god
Ordning
och
skick
tjänande
/
här
efter
framgent
behållas
/
och
ingen
ha
makt
,
av
egen
godtycke
/
däruti
något
att
förändra
;
Där
uppå
Biskoparna
och
Superintendenterna
med
DomKapitlen
,
måste
flitigt
inseende
ha
/
och
så
laga
/
att
i
alla
Stift
blir
hållen
en
Likhet
.

Texten
skall
ordentligt
/
dock
korteligen
och
enfaldeligen
förklaras
/
efter
dess
egentliga
Mening
/
med
allvarsamma
undervisningar
och
förmaningar
/
lämpade
tiIl
åhörarnas
Förstånd
/
Tröst
och
uppbyggelse
/
så
att
alla
/
enkannerligen
de
Unge
och
Enfaldige
/
må
det
grundligen
fatta
/
begripa
/
och
sig
till
förkovring
i
lära
och
leverne
/
nytteligen
anlägga
.

De
skola
vänja
sig
/
till
att
tala
rätt
Svenska
/
och
bruka
Ord
som
alla
kunniga
är
;
Och
där
de
något
i
Predikningarna
på
Latin
indraga
/
som
sällan
ske
måste
/
skall
sådant
strax
uttolkas
.

Då
skall
Gudstjänsten
börjas
med
en
morgon
Psalm
och
O
Gud
vi
lovar
dig
.

Uti
de
Vecko
Predikningar
som
ske
i
Städerna
/
skola
Texter
av
gamla
och
Nya
Testamentets
Skrifter
/
korteligen
och
grundligen
förklaras
;
Ett
helt
eller
halvt
Kapitel
åtminstone
/
som
det
är
långt
till
/
skall
uppläsas
och
uttydas
var
gång
/
och
den
Bok
som
begynnes
/
skall
ordentligt
till
ända
föras
.

Til
thessa
Veckopredikningar
i
Städerna
/
rings
första
gången
/
om
Morgonen
Klockan
sex
och
sedan
andra
gången
halvgånget
till
sju
.

Om
någon
Helgdag
infaller
på
Mån
eller
Tisdagen
/
då
blir
allenast
Bön
om
Onsdagen
;
Infaller
han
på
Torsdag
eller
Lördagen
/
sker
Bön
om
Fredagen
.

I
Städerna
hålls
då
tre
Predikningar
/
även
som
på
de
stora
allmänna
Bönedagarna
;
I
de
två
första
/
skall
handlas
om
Christi
Lidande
och
Korsfästning
;
Men
i
Aftonsången
om
dess
Begravning
.

Så
framt
uti
sättet
till
att
förrätta
Gudstjänsten
/
antingen
uti
Bönerna
/
Texterna
och
Sången
/
eller
och
själva
Tiden
/
på
vilken
Predikan
bör
hållas
/
Catechismus
förklaras
/
och
Folket
där
uti
förhöras
/
något
av
ens
eller
annans
godtycke
/
finnes
vara
för
detta
infört
/
som
intet
kommer
överens
med
denne
/
så
och
den
uti
Handboken
föreskrivna
Ordning
/
det
skola
Biskoparna
vid
Visitationer
,
och
Kyrkoherdarna
var
å
sin
Ort
avskaffa
/
samt
Allmogen
behörigen
undervisa
/
om
den
nyttan
/
som
en
likformighet
i
Gudstjänstens
övning
med
sig
har
;
brukandes
här
vid
varsamhet
och
lämpa
/
så
att
ingen
må
där
över
förargas
.

Men
på
Landet
/
skall
Folket
om
en
Söndags
Högtids
eller
stor
Böndags
Morgon
skriftas
/
sedan
Catechismi
förhör
är
förbi
/
och
förr
än
det
sammanrings
till
Högpredikan
;
Vilket
även
väl
dem
/
som
i
Städerna
boendes
är
/
skall
efterlåtas
/
om
de
det
åstunda
.

§
.
V
.
Vid
uppenbara
skriftemål
/
skall
Prästen
varna
Folket
/
att
icke
vara
så
obetänkt
/
och
förvita
den
botfärdige
Syndaren
/
det
han
Kyrkoplikt
utstått
/
och
sig
således
för
Gud
ödmjukat
har
;
Gör
det
någon
/
skall
han
därför
tillbörligen
näpsas
/
och
av
världslig
Rätt
/
med
Straff
beläggas
.

På
Stora
Högtids
Dagar
/
såsom
förste
Dag
Jul
/
Påsk
och
Pingst
/
må
inga
Bröllop
hållas
;
Men
om
någon
/
för
särdeles
skäl
och
Orsaker
skull
/
vill
i
Fastan
gifta
sig
/
bör
sådant
icke
vägras
/
allenast
det
sker
i
stillhet
/
och
utan
allt
Brudebång
.

När
årsloppet
så
medgiver
/
att
Dominica
VI
.

Sönes
det
någon
/
då
skall
han
/
sedan
Saken
i
Konsistoriet
varit
angiven
/
och
alla
medel
till
förlikning
försökte
/
förvisas
till
världslig
Rätt
/
och
Föräldrarna
vara
pliktiga
/
att
säga
sina
skäl
;
och
om
de
/
efter
noga
beprövande
gillas
/
äger
Sonen
Föräldrarna
åtlyda
.

Gör
det
någon
/
vara
sådant
ogillt
/
och
plikta
för
Brott
sin
.

Samma
Lag
var
med
de
Trolovningar
/
som
ske
med
någon
/
som
mycket
drucken
är
/
och
det
sedan
ångrar
.

Ingen
Brudskara
må
komma
till
Kyrkan
/
med
Trummor
/
skjutande
/
och
varjehanda
otjänligt
Buller
;
Sker
det
/
då
skola
sådana
plikta
efter
Stadgan
.

Om
Skillnad
i
Trolovningar
och
Äktenskap
.

Till
yttermera
visso
/
har
Vi
detta
med
egen
Hand
underskrivit
/
och
Vårt
Kungl.
Sekret
bekräfta
låtit
.

Var
alltid
redebogne
till
att
svara
varje
och
en
som
begär
skäl
etc.
Ty
vare
ock
då
denna
efterföljande
korteliga
vår
svar
i
saken
till
båda
parterna
.
,
Först
det
vi
Svenska
har
(
såsom
ock
det
samma
uti
många
andra
Kristen
land
och
Furstendöme
skett
är
)
i
många
stycken
trätt
ifrån
den
Romerska
kyrkans
stadgar
och
Ceremonier
,
är
ingalunda
skett
av
förvetenhet
,
Utan
i
sanningen
har
det
varit
oss
av
nöden
,
Ty
så
har
det
sig
med
de
Påvskas
kyrkostadgar
,
Dekret
och
Dekretal
,
så
fjärran
är
de
till
en
ganska
stor
part
,
komna
ifrån
den
enfaldighet
.
som
är
i
Christo
,
att
hon
som
helst
ha
och
behålla
vill
den
rätta
och
rena
Evangeliska
Läran
,
han
måste
sådana
stadgar
lika
som
hinderliga
och
förargliga
i
saken
förkasta
och
bortlägga
.

Här
till
skall
man
ock
räkna
de
sätt
,
Formler
och
ordningar
,
som
man
behöver
till
så
margahanda
Kristliga
handlingar
uti
Församlingarna
,
nämligen
,
till
Predikan
,
Döpelsen
,
HERrens
Nattvard
,
till
att
handla
med
de
sjuka
,
begrava
de
döda
,
skrifta
de
botfärdiga
,
bannlysa
de
tredska
och
obotfärdiga
,
Kyrkotjänare
ordinera
,
äktafolk
sammangiva
,
och
(
där
så
ske
måste
)
åtskilja
,
Ty
där
man
uti
en
Kristlig
församling
slika
vissa
ordningar
,
som
uti
våra
Agende
böcker
,
dem
vi
kallar
Handböcker
författade
är
,
icke
hade
sig
efterrätta
,
så
att
var
och
en
för
den
skull
dessa
stycken
måste
så
förhandla
,
som
honom
själv
täckes
,
eller
såsom
det
kunde
efter
lägenheten
råka
sig
för
honom
falla
,
kan
var
och
en
väl
tänka
,
vad
där
av
ville
komma
för
en
oskicklighet
,
och
församlingarna
emellan
för
en
oenighet
och
tvist
.

Icke
kunna
heller
denna
belätes
fiender
av
Skrifterna
annat
bevisa
,
än
att
beläte
icke
är
tillbedjandes
såsom
Gudar
,
efter
Hedniska
villor
,
Ty
eljest
är
själva
Skriften
full
med
beläte
,
Eller
vad
annat
är
alla
Leuitiska
Ceremonier
,
än
belätes
slag
,
genom
vilken
den
Helige
Ande
har
oss
avmålat
det
tillkommande
goda
i
Christo
?

Och
åter
en
god
tid
där
efter
,
lät
Konung
Stenkil
kalla
här
in
i
Riket
Predikare
,
synnerliga
de
två
Adelward
och
Staphan
.

Men
snälle
i
det
att
de
kunna
se
och
veta
tid
,
rum
och
andra
lägenheter
till
att
både
tala
och
tiga
,
Ty
säger
och
Salomon
,
Att
ett
ord
talat
i
rätt
tid
,
är
lika
som
ett
guldäpple
författat
i
silver
smide
.

Såsom
där
man
ville
tala
för
enfaldigt
folk
om
människornas
rättfärdighet
,
och
sade
,
Att
den
som
tror
på
Christum
,
han
är
rättferdig
,
intet
mer
tilläggandes
.

Ja
efter
menige
man
mestadels
är
så
till
sinnes
,
att
de
mer
rätta
sig
efter
gärningarna
,
som
är
för
ögonen
,
än
efter
orden
,
som
de
höra
,
skaffar
den
hos
dem
en
ringa
frukt
,
han
må
predika
så
väl
han
kan
,
som
otillbörliga
lever
,
och
således
synes
själv
ogilla
det
han
lär
,
Där
till
med
,
efter
Gud
ock
så
bär
styggelse
vid
alla
ogudaktiga
,
kan
man
icke
heller
förmoda
hans
nåd
och
välsignelse
till
den
predikan
som
en
ogudaktig
Predikare
framför
.

Och
skall
man
detta
så
förstå
,
att
innan
en
timma
skall
det
allt
ändas
,
som
en
tid
till
talande
är
,
både
förmaningen
till
bönen
,
förr
och
efter
predikan
,
så
ock
själva
predikaren
eller
utläggningen
,
eljest
var
man
gör
förmycket
långt
,
så
att
folket
begynner
ledas
vid
,
följer
där
föga
frukt
med
.

Och
förmanar
Predikaren
tillförne
folket
till
att
bedja
vid
detta
eller
något
annat
sätt
,
korteliga
.

Sedan
bett
är
,
rättar
församlingen
sig
upp
igen
,
och
står
stilla
så
länge
Lesten
eller
Texten
som
förhandlas
skall
,
är
uppläsen
.

Item
vissa
tider
,
nämligen
,
Påsk
,
och
Pingst
dagar
,
vissa
böner
,
besvärjelse
,
Evangelium
etc.
Vilket
allt
efter
det
är
fritt
och
vilkorliga
,
och
icke
hör
till
Döpelsens
rätta
väsende
,
som
uti
inga
andra
står
,
än
i
dess
egen
Ord
,
Watnena
och
Andanom
,
kunde
slikt
icke
vara
för
andra
saker
skull
gjort
,
än
att
man
således
ville
pryda
detta
Sakramentet
.

Dock
skola
samma
Barnamorskor
alltid
giva
kvinnorna
ett
gott
hopp
till
livs
,
och
icke
förfara
dem
i
deras
vånda
,
med
någon
otida
ord
om
döden
,
med
mindre
farligheten
kunde
vara
desto
större
,
Ty
när
så
är
fatt
,
då
må
de
väl
,
ja
de
måste
då
röra
där
om
,
och
giva
dem
det
in
,
Att
de
aldrig
kunna
någon
tid
bättre
dö
,
än
även
nu
medan
de
stadda
är
uti
deras
rätta
kall
,
varför
de
ock
skola
vara
fullvissa
på
Guds
nåd
och
hans
saliga
Rike
,
Där
om
ock
S
.
Paulus
rör
sägandes
,
Kvinnorna
varda
saliga
genom
barnsbörden
,
om
de
blir
i
tron
etc.
Vid
samma
sättet
skola
ock
Prästerna
förmana
havande
kvinnor
,
på
det
de
må
lära
besinna
,
att
livsfrukt
är
en
besynnerlig
Guds
gåva
,
för
vilka
de
skola
honom
med
glädje
tacka
,
alltid
befallandes
samma
frukt
,
så
väl
ofödda
som
födda
,
uti
Guds
milda
händer
,
och
innerliga
bedjandes
,
att
Gud
värdigas
sig
där
om
nådeliga
vårda
låta
.

Ty
det
är
icke
alla
,
som
uti
de
svåra
syndafall
sig
själva
veta
rätt
skicka
in
för
Gud
.

Vilken
rannsakan
är
ock
en
stor
orsak
där
till
,
att
vi
denna
hemliga
Skriftemålen
,
för
de
enfaldiga
och
unga
Kristna
skola
behålla
.

När
då
någon
som
uti
en
sådana
uppenbara
last
fallen
är
,
kommer
(
såsom
plägsed
är
)
för
Kyrkodörren
,
skall
Kyrkotjänaren
,
den
som
plägar
kallas
Pänitentiarius
,
granneliga
rannsaka
om
det
fallet
.

Item
man
må
och
väl
sätta
dem
allmosegåva
och
andra
misskundsamliga
gärningar
,
varje
som
hans
lägenhet
och
ämne
tillsäger
.

Ty
så
säger
HERren
,
Jag
ser
till
den
elände
,
och
till
den
som
har
en
förkrossat
anda
,
och
fruktar
mitt
ord
.

På
Landsbygderna
må
väl
Mässan
alltid
och
alltsammans
hållas
på
Svenska
.

Men
på
det
man
skall
icke
synas
vilja
platt
förakta
det
Latinska
tungomålet
,
eller
låta
det
platt
falla
,
vilket
dock
alla
Klerker
behöva
och
kunna
måste
,
må
ock
så
några
Latinska
sånger
,
så
väl
i
Mässorna
som
i
andra
Tider
,
brukade
varda
,
besynnerliga
i
Städerna
där
Scolar
är
,
på
stora
Högtids
dagar
eller
Apostla
dagar
.

Men
med
Mässorna
rättar
han
sig
eljest
efter
det
sätt
och
ordning
,
som
den
Svenska
Mässboken
utvisar
.

﻿För
Erick
Mickilsson
och
Per
Suensson
i
Sickelsnäs
blev
således
förlikta
och
förenade
om
någon
ägor
de
hade
till
att
träta
om
,
att
Per
Suensson
skulle
utlägga
till
allmänning
allt
vad
östen
till
vägen
var
av
en
hage
,
han
på
allmännings
mark
hade
intagit
,
det
han
och
här
på
tinget
utlovade
sig
göra
ville
.

Och
förpliktade
här
på
härads
tinget
i
nämndens
och
menige
mäns
åhöro
,
att
han
nu
strax
oförsumligen
med
hast
ville
draga
till
Stockholm
och
förskaffa
sig
sannfärdiga
brev
och
bevis
,
att
han
lagligen
hade
sig
med
sin
förra
hustru
,
för
hennes
brist
och
förseelse
som
förbe:
är
,
avskilt
.

Ändå
var
Per
Börjesson
i
Gettinge
fullmyndig
på
alla
denne
efterskrivna
syskons
vägnar
,
nämligen
:

Suen
Amundssons
i
Kulleboda
i
Lanneskeda
socken
,
Jngebor
Amundsdåtters
vägnar
i
Biedesiö
och
på
Jngridis
och
Kirstin
Amundsdöttrars
vägnar
ibidem
och
på
Heliga
och
Luze
Amundsdöttrars
vägnar
i
Glömsiö
i
Neffuelsiö
socken
och
på
Marriet
Amundsdåtters
vägnar
i
Trijshilt
i
Lanneskeda
socken
.

Kom
för
rätta
Nils
i
Byastadh
,
vilken
vart
överbetygat
,
att
han
i
förbud
hade
skjutit
en
hjort
,
till
vilket
han
icke
neka
kunde
.

Kom
för
rätta
Måns
i
Byastadh
,
som
på
nästa
framlidna
ting
utfäste
en
12
månne
ed
,
att
göra
sig
fri
för
djurskytteri
,
den
han
icke
orkade
gå
,
och
där
med
vart
han
sakfälld
till
sina
20
marker
kronan
och
häradshövdingen
till
att
böta
.

For:ne
Anna
Persdotter
hade
ingen
fångman
till
det
lärft
,
som
blev
stulet
ifrån
för:
Birge
och
blev
funnet
hos
henne
,
därmed
vart
hon
sakfälld
kronan
3
marker
och
härradshövdingen
3
marker
att
böta
.

Per
Jönsson
i
Yxeshult
Boo
i
Kärffuagårdh
Peer
i
Stocks
bärgh
Gumme
i
Lijda
Sigfridh
i
Suensholm
Måns
i
Skruff
.
hade
till
honom
,
att
han
skulle
varit
i
råd
med
en
kone
,
lille
Anna
benämnt
,
några
penningar
för
honom
att
försnilla
.

Därmed
sades
han
för
samma
tillvitelse
fri
med
mindre
någon
honom
det
skäligen
överbetyga
kan
.

Lagbudna
gårdar
Röslijda
i
Skeda
socken
2
°
Ränneridh
i
Neffuelsiö
socken
2
°
Knipshult
i
Carlstårpe
socken
2
°
Östrarp
i
Näsby
socken
2
°
Öster
gården
i
Hälleridh
i
Skeda
socken
2
°
Nörre
Knixhult
i
Kårsbärga
socken
3
°
en
fjärding
av
söndra
gården
Biedesiö
3
°
Brende
Öshult
i
Alzeda
socken
i
°
Emmeltetårp
i
samma
socken
1
°
Solshister
i
Skeda
socken
i
°
Flohult
i
Kårsberga
socken
2
°
Yxeshult
i
samma
socken
2
°
Stocketårp
i
samma
socken
30
Ekeridh
i
Huetlanda
socken
i
°
en
sättingsgård
i
Gunnarshult
i
Myresiö
socken
i
°
ANNO
1603
Den
23
juni
stod
laga
häradsting
i
Hökåsa
i
Bexeda
socken
i
närvaro
välbördig
Peer
Nilssons
till
Kulleboda
,
welb:
Nils
Jönssons
till
Åckershult
,
välförståndig
Linnert
Jörenssons
i
Hundestadh
,
kronans
befallningsman
här
i
Österhärrat
,
välaktig
Suen
Månssons
i
Rösa
underfogdes
,
hederlige
och
vällärde
mäns
herr
Ericks
i
Myresiö
och
herr
Nilses
i
Kättistårp
.

Där
om
herr
Hemmingh
allsintet
lät
sig
vårda
utan
sade
att
han
här
om
sig
ville
betänka
.

Då
kom
fram
Nils
skräddare
i
Näsby
och
gav
till
känna
,
att
fru
Beata
och
lille
Anna
skulle
ha
några
penningar
till
Näsby
och
begärde
att
hustru
Jngridh
skulle
dem
förvara
.

Detta
togs
till
rannsakning
och
bevisades
att
han
har
slagit
henne
tu
blånad
,
och
blev
för
svart
blånad
fälld
till
3
mark
.

Dock
till
det
sämste
gick
de
till
en
förlikning
så
att
de
skulle
giva
dem
ännu
oxar
3
,
var
oxe
så
god
som
4
daler
och
ett
lispund
koppar
,
och
för:ne
Måns
Gummeson
en
silversked
om
3
lod
och
hans
syster
Gunnill
Gummedoter
en
silver
sked
om
3
lod
,
här
uppå
räckte
de
händer
,
att
det
skall
vara
en
förlikt
sak
och
aldrig
här
efter
skall
påtalas
.

Nu
orsakade
samme
Jngier
sin
värbroder
Nils
Käbbeson
,
att
han
henne
aldrig
lägrat
hade
,
som
ryktet
om
honom
var
utspritt
.

Desslikes
var
Jon
i
Knixhult
fullmyndig
på
Oluffs
hustru
vägnar
i
Kiörkietårp
i
Solbärga
socken
,
att
tingsköta
Hemmingh
i
Bockebärgh
en
tolvting
av
allan
Bocke
berg
gård
för
silver
och
penningar
10
daler
.

Jtem
fram
kom
Per
Gummeson
i
Bischopsquarn
och
hans
medarvingar
och
talade
till
Jon
Alle
i
Hiupinge
torp
om
sin
broder
Jnge
Gummeson
i
Långaridh
,
som
slagen
blev
uti
et
bröllop
i
en
gård
benämnt
Engh
.

Siffridh
i
Korperydh
Gumme
i
Dale
Nils
Hemmingson
ibidem
Påffual
i
Häsleås
,
fru
en
änka
benämnt
Marriet
Suens
dotter
i
Bäxeda
och
rått
henne
med
barn
,
till
vilket
han
icke
neka
kunde
,
därför
han
vart
sakfälld
till
att
böta
kronan
,
häradshövdingen
och
häradet
penningar
2
daler
.

Därför
han
blev
sakfälld
till
att
böta
kronan
penningar
3
daler
,
häradshövdingen
och
häradet
3
daler
.

Svaranden
Item
här
uppå
utav
svaranden
befann
mann
slätt
ingen
gensvar
,
för
vad
orsaks
tillfälle
denne
förnämnde
gård
Nässiö
är
kommen
ifrån
skatten
och
skriven
in
under
kronan
,
utan
detta
ställdes
in
till
gud
,
höge
överheten
och
kammar
råd
med
kamrererna
till
att
efter
rannsaka
uti
kronans
jordlängder
.

Blev
för
det
således
interlocutorie
avsagt
,
att
Påvel
Gruvfogde
,
vilken
bemälde
Eng
för
hans
lön
gives
för
-
80
daler
kopparmynt
skall
bemälde
hö
emot
taga
,
så
mycket
han
kan
någorledes
komma
till
väga
utan
sin
Märklig
skada
antaga
,
och
Nämningeman
skall
veta
besked
på
dem
som
det
höet
bärgade
,
vilket
Påvell
sig
till
betalning
anammat
.

Vad
den
rannsakning
anlangar
,
som
Anderssboerne
därpå
hållit
har
,
och
kalla
det
en
dom
,
därefter
de
halva
mossen
slagit
hade
:
så
var
den
samma
Syn
intet
Lagligen
Nämnd
,
utan
eljest
extraordinarie
hade
befallningsman
befallit
några
av
Nämnden
där
om
rannsaka
,
vad
skäl
Parterna
ha
kunna
som
var
Rå
&
och
intet
döma
,
ej
heller
bekände
Nämnden
sig
dömt
ha
,
utan
sagt
sig
kunna
bestå
det
de
sett
har
,
och
därefter
har
Anderssboerne
slagit
till
halva
mossen
menandes
det
vara
dom
som
sagt
är
/
:
ubi
processus
nullus
,
ibi
sententia
nulla
:
/
och
det
av
missförstånd
,
och
vad
därför
för
straff
och
pen
följa
vill
,
varda
de
förnimmandes
när
om
Rågången
efter
deras
begäran
som
bemält
är
synt
och
Prövat
varder
.
10
.

besvärade
sig
accusando
bemälde
Olof
Andersson
utöver
Herr
Nillss
i
Eedboo
kyrkoherde
,
vilken
hade
handlat
med
Olofz
broder
Mårthen
om
en
oxe
,
som
sades
vara
sex
år
gammal
,
och
givit
honom
intet
mera
än
-
4
tunnor
Säd
där
dock
oxen
hörde
/
:
som
han
föregav
:
/
bemälde
Olof
till
:
begärandes
i
detta
sinne
sentens
och
Dom
:

Nu
är
omsider
så
vida
med
Saken
kommit
,
att
Härads
Syn
är
på
bemälde
ort
och
kvarnar
beviljat
och
Hållen
,
som
skedde
den
8
Juli
sist
förlden
,
uti
bemälde
stridige
Parternas
Närvaro
,
vilken
Syn
att
bevista
och
utföra
jag
undertecknat
jämte
Härads
Nämnd
25
.
extra
ordinem
befallt
var
,
ändock
jag
med
härads
hövdings
dom
havandes
Ämbets
utförande
då
här
i
häredet
intet
hade
att
beställa
.

Sedan
uppvisade
först
bemälde
käranden
,
och
sedan
svaranden
var
sin
förmente
Rågång
,
emellan
Såtter
och
Bännebool
,
men
på
ingendera
sidan
fanns
någon
Råsteen
som
vitsord
givas
kunde
,
utan
vore
ovalda
Skogsstenar
,
vad
den
Rå
anbelangar
som
stod
på
en
holme
vid
Sjöstranden
,
och
tillförne
Laggill
varit
har
,
den
vore
nu
ifrån
sitt
rätta
Rum
bortkastat
,
vilken
om
han
oförvanskat
stått
hade
,
har
han
god
Rättelse
uti
Saken
gjort
:
varför
har
Bureus
så
vitt
denna
Saken
drivit
emot
Bäncht
i
Bännebol
,
att
han
Lagfäst
har
för
samma
Råstens
uppkastande
,
den
han
ej
gått
har
.

Dirich
Keijser
som
den
tiden
skrivare
var
vid
bruket
,
bekände
sig
bemälde
tionde
av
Mårthen
ha
bekommit
,
dock
ville
han
det
intet
Befallningsman
gottgöra
förra
än
han
får
kvittensen
igen
,
som
alldeles
förfaren
är
,
antingen
av
befallningsman
eller
Mårthen
,
Blev
omsider
avsagt
,
att
medan
Dirich
Keijser
bekände
sig
Spannmålen
ha
bekommit
,
blev
befallningsmans
tilltal
på
Nämningeman
kraftlöst
,
eljest
skedde
honom
förnär
,
om
han
Säden
andra
resan
betala
skulle
,
efter
Dirich
Keijserss
Protestation
:
jämväl
erkändes
Keiser
bemälde
Spannmål
befallningsman
avhöra
,
oansett
kvittenset
är
förkommet
.

Och
efter
Olof
intet
kunde
efter
betänkande
värjas
,
erkändes
han
med
Laga
Ed
sig
och
sina
befria
,
att
de
icke
vore
orsaken
till
hästens
fördärv
,
när
det
skett
är
,
varder
Saken
emot
knekten
om
han
lever
,
utförd
.
33
.

besvärade
sig
klageligen
bemälde
Madz
Erichsson
över
bemälde
Peer
Staphansson
som
honom
för
tjuveri
beryktat
hade
som
förra
akta
utvisa
,
Peer
svarade
sig
beskyllningen
kunna
bestå
och
vilja
bevisa
honom
sina
Kattiskor
stulit
ha
,
vilket
när
han
med
vittnen
försöka
skulle
,
nekade
de
icke
allenast
till
det
Per
dem
om
samma
tillmäle
åtsporde
sig
till
hjälp
reda
,
utan
bekände
offentligen
sig
intet
annat
veta
med
bemälde
Madz
Erichsson
än
det
som
ärligt
var
;
och
efter
såsom
bemälde
Per
Staphansson
sig
ej
rätta
ville
,
utan
beskyllningen
påstod
,
och
det
ej
bevisa
kunde
Sakfälldes
han
till
-
40
₥
Tingmale
B
:

kom
för
Rätten
Thomass
Andersson
i
Järssöö
uti
Kasskyrkie
Socken
,
och
på
välborna
Fru
Brijta
Bielkess
etc.
vägnar
kärade
till
välbetrodda
Fru
Jngeborgh
Ulfsparress
etc.
mjölnare
.

berättade
Nämnden
sig
jämte
underLagmannen
välaktat
Olof
Mårthensson
,
ha
varit
kallade
till
Gufvesta
där
till
åtskilja
några
tvistigheter
,
som
emellan
Larss
Cnutzson
och
Madz
Grijss
svävat
har
,
angående
en
slåtthage
,
vilken
Larss
Cnutzson
nu
klandrar
och
förmenar
att
Kronohemmanet
där
han
bor
skall
vara
något
preiudierat
,
och
dömt
att
Kronohemmanet
där
Larss
bor
har
sin
fullnad
emot
bemälse
hage
annorstädes
.

kom
för
Rätten
Erich
Thomasson
vid
Orthale
och
klagade
till
hustru
Charin
i
Lingslätt
,
som
hade
med
en
häst
kört
på
hans
moder
hustru
Elin
,
att
hon
föll
vid
isen
,
och
därför
en
tid
hållit
vid
Sängen
.

Och
medan
sådana
granne
trätor
pläga
ofta
stor
vidlyftighet
förorsaka
,
sattes
vite
dem
emellan
vid
-
40
₥
,
sådant
i
tid
att
avskaffa
och
förhindra
.

Och
vidare
skall
rannsakas
om
de
några
Svedjeland
huggit
har
och
där
några
Ekar
antingen
fällt
eller
och
förbränt
genom
försummelse
eller
eljest
bevåg
,
när
det
skett
är
varder
Dom
ågiven
.
etc.
55
.

Tre
drängar
i
VästerNääss
Sakfälldes
till
3
₥
för
svarslösa
stämda
för
tjuveri
på
Rovor
etc.
S
:
D
:

gav
Madz
Mjölnare
vid
Järssiö
tillkänna
sig
ha
vederkänts
hos
hustru
Brijta
i
Össbytorpedt
,
en
Skinkassjacka
,
och
en
vallmarsströja
,
vilka
för
sex
år
sedan
ibland
mycket
annat
honom
ifrånstulna
blev
,
vilka
hon
bekände
sig
köpt
ha
,
och
den
dem
sålde
,
bekände
Madz
intet
vara
sanna
tjuvar
.
hos
honom
som
henne
dessa
persedlar
sålt
har
skall
vidare
erfaras
och
Rannsakas
,
hur
han
sådant
bekommit
har
,
och
om
den
kan
därigenom
uppsynas
som
honom
stulit
har
;
och
föregivs
den
bo
uti
Väddöö
Socken
,
som
skall
vara
hennes
fångeman
.
77
.

kom
för
Rätten
manhaftig
Per
Larssonss
i
Nääss
uti
Bro
Socken
,
fullmäktig
för
Jonas
Khönichsson
,
och
begärde
av
härads
Nämnd
Dom
på
den
Lagkallade
Synen
,
som
den
10
Maj
hållen
blev
,
emellan
bemälde
Löjtnant
och
hans
grannar
Anderss
Madzson
samt
Erich
Larsson
,
alla
kärande
.
och
Ekebyborna
samtliga
svarande
,
anlangande
en
Ström
vid
utgrunds
Bron
,
som
Ekebyborna
här
till
innehaft
och
brukat
har
.
där
dock
Nässbornas
ägor
och
Äng
är
på
den
ena
sidan
om
Saxvijken
och
Strömmen
emot
bemälde
Ekeby
.

Nämligen
att
enär
bemälde
Marcus
var
i
ett
gästbod
i
Gåfvesta
,
hade
han
om
en
Natt
besovit
bemälde
Chierstin
i
bagarstugan
i
Högsätet
,
ty
hon
Låg
där
förre
,
och
när
han
inkom
gick
han
strax
dit
;
då
tillspordes
denne
Olof
,
om
han
sådant
varse
blev
,
eller
vilken
mera
då
i
stugan
var
,
han
svarade
att
folket
sov
,
men
en
hustru
,
benämnd
Margaretha
satt
i
spisen
,
och
vet
grant
här
om
sade
han
berätta
;
vidare
fann
han
dem
intet
i
gärningen
,
än
att
han
hörde
Marcus
Spårar
ringa
som
en
klocka
;
Till
detta
Nekade
både
Han
Såsom
och
denne
Chierstin
.

Mera
att
bekänna
kunde
han
honom
intet
övertala
eller
beveka
,
Nu
tillspordes
han
,
vad
han
här
till
svara
ville
;
han
gav
det
svaret
ifrån
sig
,
att
han
allenast
tänkte
denne
lede
gärningen
göra
,
och
var
han
hade
icke
blivit
förhindrat
,
likväl
fullborda
.
på
detta
stod
han
allt
stadigt
.

Då
blev
Predikanten
uti
Rassboo
förordnat
honom
ensligen
förmana
till
sanningens
bekännelse
,
då
kom
han
omsider
så
vida
med
honom
,
att
han
sade
sig
och
före
ha
haft
i
sinnet
sådant
bedriva
med
ett
Sto
hos
sin
husbonde
Anderss
Olofzson
,
och
intet
vidare
det
fullföljt
,
eller
så
när
kommit
som
med
bemälde
andra
Kreatur
.

Sedan
åter
in
för
Rätten
bekände
han
efter
foglig
föregången
förmaning
,
att
han
tre
resor
sig
med
Stoet
uti
sin
Matfaders
Stall
beblandat
har
Näst
för
sista
våren
,
och
att
ingen
hade
det
varse
blivit
,
men
med
det
andra
Kreatur
,
intet
mera
än
den
ena
resan
dock
fullkomligen
etc.
mera
eller
med
flera
Kreatur
bekände
han
intet
,
ej
heller
blev
honom
sådant
övertygat
,
mycket
mindre
hade
där
till
honom
någon
tubbat
.

Såsom
ock
den
Högstberömligaste
Kungl:
Hovrättens
i
Stockholm
av
gångne
brev
Dat
:
6
Maj
om
den
Unge
Skrivaren
\
Hans
Johansson
/
som
har
ihjäl
slagit
Överstelöjtnanten
Erich
Reuter
,
att
den
honom
kunde
fast
bringa
,
skall
bekomma
en
ansenlig
penning
summa
.

Hindrich
begär
och
där
hos
av
Sannfärdigt
Skottsmål
och
vittnesbörd
om
sitt
före
hållande
den
tid
han
här
i
Socknen
varit
har
,
vilket
där
och
alla
vedermän
gjorde
,
att
han
sig
hos
dem
tro
ärligen
och
redligen
förhållit
har
den
tid
han
hos
dem
vistas
har
Såsom
och
framtändes
ett
vittnes
börd
,
av
be:te
Spores
broder
honom
givit
den
han
tjänat
har
uti
en
tid
,
att
han
honom
troligen
tjänat
har
,
och
icke
vet
heller
kan
honom
i
några
måtto
att
beskylla
hel:r
beklaga
.

Och
Siul
och
Erich
Olufssönner
skola
igen
lägga
de
6
.
orter
som
de
utav
honom
på
Köp
uppburit
har
,
helst
efter
de
icke
kunna
frälsa
eller
hemula
honom
på
hela
gården
.

Upplästes
Kungl.
Maij:tz
Drottning
Christinæ
Resolution
och
förklaring
à
Dato
Stockholm
d
.
27
Februari
A:o
1653
angående
alla
Pantgods
Reduktion
,
till
dess
rätta
odel
eller
Bolbyer
.

Blev
om
Jon
Olofsson
i
Biörsiö
Käromål
om
...
Hemmanets
inlösande
slutit
,
att
efter
han
störste
delen
av
Samme
Hemman
inlöst
haf:r
behåll
...

(
17
.
)
Uppbjuder
Nilss
Ifwarsson
i
Bågsiö
andha
gången
Slåttänget
Östbyn
för
14
RikD:r
inlöst
.

Cap.Landzl:n
så
och
Hans
Höggrefl:e
Excell:tz
H:r
Guvernörens
Högvälborne
H:r
Carl
Sparres
givna
instruktion
,
Daterat
Sunne
den
3
Maj
A:o
1666
.

Erik
Pehrson
i
Flattnohr
Anderss
Olufson
i
Grönuiken
Tohl
Nillson
i
Sidsiöö
Pehr
Bengtson
i
Biörnöhn
Nillss
Nillson
i
Molvuiken
Brodde
Olufson
i
Rindh
.

Biörnöhen
skall
därför
plikta
3
mk:r
Sm:tt
för
vartdera
efter
33
Kap
Tingb:n
LL
.

Efterskrivna
Bräcke
bor
som
ej
haf:r
avlagt
sin
fiske
tionde
hos
kyrkoherden
,
utan
än
restera
,
såsom
Nillss
Nillsson
i
Mohlwijken
för
6
år
,
Oluf
Michelsson
för
7
år
,
Oluf
i
Bröcklinge
för
8
år
,
Månss
Olufsson
i
Beensiö
för
4
år
,
Erich
Erichsson
ibid
.
för
6
år
,
Anders
Olufsson
för
4
år
,
men
tillstår
allenast
ett
år
,
de
övriga
inständigt
nekar
till
emot
kyrkoherdens
tionde
Längds
bok
,
Oluf
Carlsson
för
7
år
,
skulle
var
om
sig
plikta
för
treska
och
emot
vilja
var
sina
3
mk:r
S:m:tt
belöper
21
mk:r
och
Månss
Olufsson
för
flärd
3
mk:r
för
oduglig
upprutten
fisk
var
med
de
för
denne
gången
förskonades
.

Länsman
Pehr
Andersson
betygade
med
själv
sina
eder
att
han
till
sal
.

Anno
1673
den
10
Oktober
,
Hölls
Laga
Ting
i
Rääfsundz
Giäldh
,
Närvarandes
Kronans
Befallningsman
Wälb:de
Daniel
Bertilsson
,
tillika
med
de
Tolv
Edsvurna
Nämndemän
.

Johan
Trumslagare
betygar
och
,
om
13:de
dags
Morgon
då
han
inkom
i
Storstugan
,
stod
Kapten
Anrepp
och
tvättade
sig
,
sade
han
,
skulle
en
sådan
Hundzfott
föra
sina
Horor
in
på
mig
.

Förelästes
Tolvmäns
Rannsakningen
emellan
Kyrkoherden
Vördig
och
vällärde
H:r
Isaac
Alstadium
och
hans
Son
H:r
Carl
,
å
den
ena
sidan
Kärande
och
Kapten
wälb:
Gosvin
Anrepp
å
den
andra
Svarande
,
som
hållen
blev
den
10
Oktober
1673
Vilken
Rannsakning
Tolvmän
,
ord
ifrån
ord
vederkände
,
så
vara
passerat
,
som
i
Rannsakningen
annoterat
och
infattat
är
,
och
icke
förstå
kunna
till
det
ringesta
något
vara
förgätit
,
Vilket
de
med
Ed
erhålla
vilja
,
när
så
fordras
,
Fördenskull
de
sitt
Gäldens
Signet
samtyckte
samma
Rannsakning
att
verifiera

Pehr
Olufsson
i
Noor
klagade
,
huruledes
Fogdekarlen
Lars
Falk
har
några
veckor
för
Påsk
illa
slagit
och
hanterat
sig
,
när
han
kom
körandes
ifrån
Noor
och
till
Döfwinge
,
ämnandes
köra
till
Bådsiö
efter
Råg
,
när
han
om
afton
sent
inkom
till
Döfwinge
,
som
var
hans
Fars
gård
,
att
begära
hus
,
vore
där
för
honom
Länsman
Pehr
Andersson
och
Lars
Falk
inne
uti
Stugan
,
då
har
Lars
Falk
begynt
ajera
honom
,
efter
han
satte
sig
fram
på
bänken
,
Lagt
hyend
fram
,
bett
sitta
när
han
har
vägrat
,
tagit
i
håret
och
slagit
,
som
Lars
Falk
här
ifrån
ej
kunde
neka
,
utan
bekänner
så
vara
skett
,
vilket
och
Länsman
Pehr
Andersson
tillstod
ha
dem
skilt
åt
,
då
har
Pehr
Olufsson
sedan
utgått
att
gömma
sig
undan
i
ett
Stall
där
Gårdshästarna
stod
,
där
inne
var
och
Lars
Falkz
Fohla
,
har
Falk
kommit
efter
löpandes
och
fann
där
åter
Pehr
Olufsson
för
sig
i
Stallet
,
strax
tagit
i
Håret
,
slagit
i
golvet
och
Spänt
på
veklivet
Lars
nekar
,
ha
honom
sparkat
,
utan
allenast
Hårdragit
och
Pustat
,
inga
vittnen
,
har
det
på
sett
,
Vad
som
i
Stallet
var
passerat
.

Oluf
Andersson
i
Mälbyn
på
Frössöön
på
Lars
Olufsons
wäg:r
ifrån
Rijse
fordran
3
RD:r
lånade
Penningar
och
1
Spann
Korn
,
av
Snickarens
sal
.

Kronans
Befallningsman
wälb:de
Jonas
Flodin
besvärade
sig
hur
\
han
/
en
och
annan
tid
har
fått
skriftliga
tilltal
av
Hans
Excell:z
Högwälb:e
H:r
Guvernören
om
Postlöpandets
oriktiga
fortgång
,
här
igenom
Räfsundz
Tingslag
,
förehölls
alltså
Pehr
Andersson
Länsman
,
som
och
Post
bonde
är
,
hur
det
till
kommer
,
varutinnan
försumnelse
sig
består
,
giver
anledning
det
Swen
Nilsson
i
Bräcke
skicka
honom
gård
emellan
ifrån
Bräcke
,
och
i
synnerhet
nu
senast
skickat
med
Gååsböhle
flickan
;
som
och
alltsomoftast
tillförne
sänt
Posten
om
Söndagsmorgon
med
Grimnäs
Kyrkfolket
till
Räfsundz
länsmansgård
.

Nills
Jonsson
i
Mälgåsen
,
Siuhl
Sedfastson
i
Tamnäs
Fast
Persson
i
Böhle
,
Bengt
Persson
i
Marset
Oluf
Persson
i
Fanbyn
,
Kiehl
Persson
i
Giällön
Herman
Person
i
Biöröen
,
Nills
Persson
i
Anwijken
Erich
Andersson
i
Ring
,
Lars
Larsson
i
Beensiö
Pehr
Andersson
i
Sidssiö
Pehr
Olsson
i
Grimnäs

(
19
)
Proviantmästaren
Peder
Erichsson
Niure
lät
uppvisa
Tvenne
sina
förlängst
lagbudna
och
lagståndna
Köpe
brev
på
Lanssom
gård
,
av
Oluf
Ersson
Ibm
på
halva
gården
och
den
andra
halva
delen
till
Kreditorerna
efter
Härads
Rättens
Resolution
d
.
5
Juni
1679
inlöst
;
Varför
beviljades
honom
på
hela
hemmanet
Dombrev
.

L.L
.
till
sig
lösa
,
det
övriga
av
Hemmanet
hör
Sonen
Jöns
Jonson
till
,
som
är
gift
i
Norie
och
Dottern
Märitt
Jonsdotter
och
Tårckell
stiger
således
där
ifrån
.

Och
de
trädde
uti
förbundet
,
att
de
skulle
söka
HERREN
,
deras
Faders
Gud
av
allt
hjärta
,
och
av
all
själ
,
Och
vilken
som
icke
sökte
HERREN
Israels
Gud
,
han
skulle
dö
,
både
liten
och
stor
,
både
man
och
kvinna
.

Och
på
det
att
samme
Religions
Bekännelse
,
må
så
väl
främmande
som
infödda
kunnig
vara
,
Därför
vart
i
själva
Konsiliet
beslutat
,
såsom
vi
ock
nu
för
nyttigt
,
nödigt
och
rådsamt
aktar
,
att
låta
förbenämnde
Kristliga
Religions
och
vårLärdoms
förening
,
samt
med
de
tre
Guds
Församlings
tros
Bekännelser
,
vilka
Symboler
kallas
,
såsom
ock
den
rätte
,
rene
och
oförändrade
Augsburgiske
Konfession
,
vilken
Anno
etc.
30
,
på
den
store
Riksdag
,
som
då
av
Chur-Furster
och
Städer
hållen
blev
,
vart
överantvardat
Kejsare
Carl
den
Femte
,
av
Trycket
låta
utgå
:

Därför
må
vi
den
i
våra
Församlingar
efter
en
Kristen
friheet
väl
bruka
.

Såsom
icke
heller
något
annat
av
de
Påskas
lärdom
eller
villfarelser
,
evad
namn
de
helst
ha
kunde
,
någon
tid
gilla
eller
vedertaga
,
utan
dem
alldeles
förkasta
,
såsom
människostadgar
,
för
världslig
höghet
,
välde
,
makt
,
och
rikedomar
upptänkta
,
igenom
vilka
många
människor
ofta
är
bedragna
vordna
.

Och
där
som
själva
saken
så
kräver
,
må
det
som
yttermera
behövs
,
med
Bisparnes
och
Kapitlens
gemena
samtycke
,
bli
tillagt
och
förmerat
.

Likväl
efter
sådant
för
handel
och
vandel
skull
icke
väl
kan
förhindrat
varda
,
så
är
så
vitt
samtyckt
,
att
dem
som
någon
Kättersk
lärdom
har
,
icke
skall
tillstått
eller
efterlåtit
vara
,
att
hålla
några
uppenbara
Samkväm
i
hus
eller
annorstädes
,
så
framt
var
några
där
med
befinns
,
eller
de
som
eljest
försmädligen
talar
om
vår
Religion
,
de
skola
tillbörligen
straffade
bli
.

Och
på
det
,
att
alla
må
kunnigt
och
veterligt
varda
,
vad
vi
ytterligare
uti
denne
Samkväm
handlat
och
oss
ha
förenat
om
,
uti
alla
Punkter
och
Artiklar
,
så
skall
sådant
med
första
av
Trycket
utgå
.

SYMBOLVM
APOSTOLICVM
JAg
tror
på
Gud
Fader
allsmäktig
,
himmelens
och
jordens
Skapare
.

Varken
sammanblanda
Personerna
,
eller
åtskilja
det
Gudomliga
väsendet
.

Item
de
som
föregiva
,
att
några
uti
detta
livet
,
kan
en
sådana
fullkomlighet
vederfaras
,
att
de
intet
synda
kunde
.

Varför
varda
ock
de
fördömda
,
som
lära
,
att
Sakramenten
göra
oss
rättfärdiga
ex
opere
operato
,
Det
är
,
allenast
för
det
omak
skuld
,
att
man
går
till
Sakramenten
,
dock
utan
tron
.

Dock
varder
folket
om
slika
stadgar
förmanade
,
att
samveten
icke
skola
bli
besvärade
,
lika
såsom
sådana
Ceremonier
vore
en
nödig
Gudstjänst
till
saligheten
.

Varför
ock
Klosterlöften
,
och
stadgar
om
åtskillig
mat
och
dagar
,
etc.
upptänkta
till
att
förtjäna
Guds
nåder
,
och
tillfyllestgöra
för
synderna
,
är
alldeles
onyttiga
,
och
motsträva
det
heliga
Evangelium
.

För
ty
,
ändock
människan
någorledes
kan
uti
utvärtes
måtto
Guds
bud
hålla
:

OSS
varder
falskeligen
tillmätt
,
att
goda
gärningar
hos
oss
förbjudna
blir
.

Vidare
varder
av
våra
Predikanter
lärt
,
att
man
måste
göra
goda
gärningar
,
icke
för
den
skull
,
att
vi
skola
förtrösta
oss
genom
dem
förtjäna
Guds
nåder
,
utan
därför
,
att
det
är
så
Guds
vilja
.

Ty
både
är
de
Konungar
.

Men
denna
sedvanan
är
icke
allenast
emot
den
heliga
Skrift
,
utan
ock
emot
Canones
eller
den
gamla
Kyrkolagen
och
Guds
Församlings
Exempel
,
i
bruk
kommen
.

Och
samme
sak
blev
sedan
så
otillbörliga
och
skamliga
handlat
,
att
icke
allenast
Äktenskap
där
efter
blev
Prästen
förbjudet
,
utan
ock
de
som
Äkta
vore
,
blev
var
ifrån
annan
skilda
,
emot
all
,
både
Guds
lag
och
mänsklig
lag
,
som
icke
allenast
av
Påvarna
,
utan
ock
av
lovvärde
Konsilj
s
och
allmänna
Möten
ärgjorda
och
stadgade
.

Så
är
icke
allenast
av
S
:

Drar
Hans
Nåd
Er
till
minnes
som
och
förmanandes
är
att
i
det
icke
förgätit
har
i
vad
punkter
Riket
och
dess
Inbyggare
uti
staden
var
/
den
tid
Hans
Nåd
kom
först
till
Regementet
/
så
att
var
Gud
icke
hade
hjälpt
och
styrkt
honom
i
det
han
företog
emot
Konungen
etc.
då
hade
icke
annan
på
färde
varit
än
alla
ers
fördärv
som
väl
på
syntes
i
den
okristliga
handel
som
K
.
etc.
här
i
landet
bedrev
med
hängande
/
brännande
/
steglande
.
etc.
till
dess
att
det
hade
väl
räckt
till
oss
alla
/
om
han
hade
längre
vid
makt
blivit
.

Och
som
h
.
N
.
sa
sig
ingen
tröst
på
färde
vara
/
annan
än
av
Gud
och
Sweriges
allmoge
den
dock
nog
försvagat
ock
förtryckt
var
av
den
stora
skada
de
lidit
hade
på
långa
Fredag
vid
Uppsala
och
i
andra
släktingar
och
där
till
med
mist
deras
armborst
och
värjor
.
etc.
Stockholm
stad
och
all
Slotten
Calmarna
/
Stägeborgh
och
tesliges
Finland
var
i
fienders
händer
/
begynte
h
.
N
.
betänka
att
Svenske
män
var
försvaga
till
det
företaget
var
och
därför
begynte
han
vinnlägga
sig
att
dra
sig
och
Riket
vänner
till
i
främmande
land
(
besynnerlig
med
Lubech
stad
och
de
andra
vendiska
städer
/
vilka
h
.
N
.
med
stort
plats
och
vedermöda
bevekade
där
till
att
de
och
trädde
in
i
saken
emot
K
.
etc.
Ty
de
vore
där
ganska
om
lwge
till
i
förstone
för
det
stora
anhang
skull
som
K
.
etc.
hade
på
Kejsarens
vägnar
/
Margreffuen
och
andra
mäktiga
Furstars
vägnar
/
dock
på
sistone
föll
de
till
h
.
N
.
och
Riket
och
skickade
här
in
skepp
/
bössor
och
värjor
/
Ryttare
och
Knektar
/
som
på
den
tid
väl
av
nöden
var
/
med
ingen
ringa
bekostnad
den
än
nu
icke
alldeles
betalad
är
.

Denna
epters:ne
framsättningar
ger
vår
nådiga
Herre
Er
Riksens
Råd
för
och
menige
Adeln
och
andra
goda
män
som
av
menige
Allmogen
här
församlade
är
i
Westras
.
etc.
Först
tackar
Hans
Nåd
Er
alla
för
Er
välvillighet
,
att
i
efter
Hans
Nåds
kallelse
komna
är
här
till
mötes
/
utan
tvivel
med
stor
kost
och
tärning
/
och
ger
er
alla
tillkänna
att
det
icke
skett
är
utav
någon
lätthet
utan
av
uppenbara
nöd
och
för
viktiga
saker
skuld
/
som
i
nu
här
skulle
få
höra
.

Och
var
han
något
mera
hade
varit
till
alders
kom
men
och
hade
vi
det
så
mycket
av
slika
landens
lägligheter
hade
han
visserligen
aldrig
givit
sina
samtycke
där
till
.

Men
h
.
N
.
höll
sig
allenast
vid
allas
Ers
löfte
/
bepliktelse
och
ed
/
som
alla
på
hela
Riksens
vägnar
h
.
N
.
där
gjorde
/
med
stor
bön
/
att
han
icke
skulle
förlåta
Er
yttermera
/
var
h
.
N
.
mesta
hop
att
Svenska
män
skulle
nu
kunna
väl
besinna
sig
av
den
vedermöda
och
obotlig
skada
och
fördärv
/
de
då
lidit
hade
/
att
de
skulle
testa
bättre
kunna
där
efter
vakta
sig
för
inbördes
tvedräkt
och
stämpling
/
och
icke
hastigt
åstunda
någon
förvandling
/
därför
för
Er
bön
skuld
och
dråpliga
bepliktelse
gav
h
.
N
.
då
på
sistone
samtycke
därtill
/
det
honom
sedan
tid
och
ofta
ångrat
har
.

Och
beklagar
h
.
N
.
sig
/
att
ändå
h
.
N
.
vinnlägger
sig
dag
och
natt
om
Riksens
bästa
/
bär
där
sorg
och
många
vaknätter
före
/
varder
dock
h
.
N
.
allt
väntan
till
det
värsta
/
så
att
där
han
förmoda
sig
tack
och
gunst
/
där
förnimmer
han
förtal
/
stämpling
och
obestånd
före
/
allra
mest
uppe
i
Dalarne
/
vilka
sig
och
berömma
att
de
har
satt
h
.
N
.
i
Högsätet
/
tackandes
sig
tillfälle
därav
att
de
var
med
när
Gud
gav
h
.
N
.
den
första
sägren
i
den
slaktning
här
i
Westrås
/
än
dock
de
gick
strax
mest
alla
hem
igen
/
och
var
då
all
Slotten
Stockholms
stad
och
allt
Finlandh
i
fiendernas
händer
/
vilka
sedan
med
menige
Riksens
tillhjälp
och
icke
med
Dalernes
allena
inkräktat
vorde
/
dock
förnimmer
h
.
N
.
att
samma
Dalakarla
mena
allt
av
deras
konst
skett
vara
/
och
att
de
för
den
skuld
vilja
och
skola
insätta
och
avsätta
i
Riksens
regemente
vem
dem
synes
/
och
därför
var
några
vill
begynna
något
obestånd
i
Riket
/
behöver
han
icke
annat
göra
än
giva
sig
upp
i
Dalarna
/
och
så
har
man
strax
uppsköt
och
nytt
regemente
/
på
vilket
ingen
lyster
vara
Riksens
Herre
/
när
han
alltid
skall
reda
sig
på
slika
vmunediga
/
och
kan
heller
då
ingen
ting
taga
sig
före
om
Riksens
bästa
/
utan
skall
alltid
vara
bekymrad
;
Om
sådana
stycken
bör
väl
övertänkas
/
om
Sweriges
Rike
skall
alltid
regera
sig
efter
dem
/
och
dem
ha
för
Herren
som
dem
av
Dalarna
uppsätter
varder
.

Har
och
samme
Dalakarle
tagit
en
sid
förre
/
att
när
en
förrädare
ger
sig
upp
till
dem
/
tager
de
honom
i
försvar
/
och
icke
vilja
låta
honom
komma
till
rätta
/
på
vilket
mången
skalk
drister
sig
ock
må
onäpst
göra
allt
det
förräderi
som
honom
lyster
/
ville
h
.
N
.
gärna
veta
/
varför
de
skola
ha
sådana
privilegier
mera
de
än
andra
lands
ändar
/
Rikena
till
så
stor
obestånd
.

Varda
desslikes
skalkar
och
stämplare
förmycket
betrodda
i
landet
enkannerliga
där
uppe
i
de
lands
ändar
/
och
må
för
den
skuld
säga
h
.
N
.
och
vem
de
vilja
allt
dem
lyster
/
det
dock
var
god
man
både
att
straffa
och
icke
lida
/
besynnerliga
medan
slika
brev
och
bepliktelse
där
om
gjorda
är
som
förberört
är
.

Så
och
för
slika
inbördes
obestånd
h
.
N
.
alltid
på
stämplas
ibland
hans
egne
allmoga
/
som
ock
nu
nyligen
skedd
är
i
Wästergötlandh
där
utsände
är
budkavla
svarade
och
brände
ibland
allmogen
/
och
har
uppropat
ett
lögnaktigt
rykte
att
h
.
N
.
har
pålagt
en
ny
beskattning
över
Riket
IIII
.

Förs
h
.
N
.
och
uppå
att
han
bryter
ned
Kyrkor
och
Kloster
det
dock
icke
finns
med
sanning
/
än
dock
väl
sanningen
är
att
Stockholms
borgare
med
stor
skäl
har
talat
om
de
Kyrkor
på
Malmarna
ligga
staden
till
stort
förfång
då
han
belagt
är
/
och
fienderna
till
godo
/
och
tyckte
intet
orätt
vara
/
att
de
nedbryts
/
vilket
dock
icke
än
nu
här
till
dags
har
varit
tillstått
.

Om
alla
föreskrivna
stycken
de
h
.
N
.
påförda
är
/
både
de
där
uppräknade
är
eller
eljest
h
.
N
.
påförs
/
är
h
.
N
.
överbödig
stå
till
svars
och
rätta
för
Er
/
och
så
reda
sig
där
ut
/
att
han
väl
hoppas
sig
försvara
i
är
och
rådlighet
/
som
en
Kristen
Furste
bör
att
göra
/
och
har
för
den
skuld
endeles
stämt
detta
möte
och
bjuder
var
och
en
som
honom
har
något
skylla
eller
till
att
tala
att
han
det
dristliga
gör
/
där
h
.
N
.
gärna
vill
tillsvara
/
med
all
rådlighet
och
Har
det
också
utskrivit
besynnerlig
upp
i
Dalarna
.

Det
väl
märkandes
att
det
icke
vill
lyckas
utan
med
allas
vår
skada
och
fördärv
/
vilket
h
.
N
.
nådigt
säger
efter
hans
av
Guds
hjälp
har
kommit
Riket
i
rolighet
och
sin
frihet
igen
/
och
ser
fördenskull
icke
gärna
att
det
skall
komma
åter
i
något
)
obestånd
igen
i
hans
tid
.

Var
för:ne
saker
icke
vår
de
h
.
N
.
enkannerliga
anröra
/
är
dock
nog
andra
saker
som
ej
allenaste
honom
utan
eehoo
han
helst
är
som
Riket
i
värjo
har
en
styggelse
skall
göra
vid
regementet
/
vilka
nu
här
efter
följa
.

Först
att
Kronans
Ränta
är
intet
så
står
som
somliga
mena
/
att
där
med
kan
hållas
så
mycket
folk
som
denne
oroliga
tider
tillkräver
/
bössor
/
värjor
/
skepp
/
harnesk
.

Kräver
och
Konungsligt
stått
mera
bekostnad
än
en
slet
Gubernatoris
,
skall
och
ofta
utskickas
sändebud
till
Herrar
och
Furstar
/
Städer
.
etc.
Och
ofta
undfångas
deras
Sändebud
igen
det
ingen
ringa
ting
kostar
/
och
sänds
nu
och
komma
desto
flera
Sändebud
och
dess
oftare
att
Riket
är
kommet
till
stadga
under
en
viss
Herre
ock
Konung
/
och
besynnerliga
då
män
vinnlägger
sig
/
(
som
h
.
N
.
nu
gjort
har
)
att
draga
sig
av
Rikena
vänner
till
med
Herrar
och
Furstar
.
etc.
Land
och
Städer
/
evar
man
kan
som
väl
nyttigt
är
.

Är
och
Slotten
förfallen
och
somliga
omkullslagen
som
för
ögon
är
där
och
ingen
ringa
kostnad
tillhör
/
om
de
uppbyggas
skulle
/
som
väl
av
nöden
är
/
både
för
inländsk
upplopp
skull
/
så
ock
för
främmande
fiender
skull
/
om
de
här
komma
.

Efter
Riddarskapet
(
som
nu
Gud
dess
lov
växer
till
igen
)
är
mycket
försvagat
för
mycket
orolig
skull
/
där
deras
gods
har
dem
avhänt
varit
med
brand
och
ville
och
mest
där
av
att
deras
gods
och
ägodelar
är
störste
delen
kommen
under
Kyrkor
/
Kloster
/
Prebender
/
begangilse
.
etc.
ville
alla
ha
hjälp
och
förläningar
)
som
intet
under
är
)
av
Kronan
och
är
då
sedan
Konungens
del
desto
mindre
till
att
upphålla
alla
för:ne
ting
.

Och
låter
h
.
N
.
er
förstå
sör:ne
stycken
inte
har
föregivit
utav
någon
lätthet
eller
för
något
snack
eller
omslag
skuld
/
utan
av
rätta
allvarliga
mening
/
att
I
må
desto
allvarligare
här
utinnan
betänkta
vara
/
h
.
N
.
känner
bäst
var
det
håller
/
h
.
N
.
tänker
och
väl
att
han
för
Riket
skuld
är
kommen
i
vilja
med
somliga
/
utländska
/
i
ty
att
han
icke
allsinget
låter
träda
på
sig
/
eller
Riket
/
skall
han
det
sedan
vänta
sig
ont
av
sina
egna
/
då
sitter
han
emellan
två
elda
/
och
gör
icke
visliga
om
han
längre
bryts
här
med
.

Munkar
som
Ränta
har
/
gick
intet
ut
att
ligga
.

Och
avläggs
den
seden
/
att
när
Prästen
dör
/
tar
Biskopen
hans
Ägodelar
/
rätta
Arvingar
till
Förfång
/
och
ger
icke
Präster
annorlunda
Testamente
/
än
efter
Lagboken
/
som
andre
Dannemän
.

Matz
Andersson
i
Hwsby
för
svarslöse
Erich
(
Bchsson
)
i
Burunge
var
vitt
av
Per
Matsson
att
han
skall
ha
tagit
honom
några
(
Rafwar
)
ifrån
Feste
lag
själv
tredje
till
näste
ting
att
göra
sig
fri
.

Vilket
ärende
jag
satte
till
Nämnden
att
rannsaka
efter
noga
rannsakan
berättades
att
då
han
vart
sack
tjänade
han
h
.
K
.
M:t
vår
Nådigaste
Konung
(
för
en
Böss
smed
därför
han
fick
lön
)
,
och
icke
(
tjänade
i
Morthen
i
Karby
)
h
.
Anna
i
Abyggeby
var
kommen
i
tal
att
hon
skulle
kunna
umgås
med
trolldom
där
om
vart
rannsakat
,
och
fanns
ingen
som
visste
av
vem
det
talet
var
utkommet
,
och
medan
ingen
var
som
kunde
henne
det
till
Lägga
,
icke
visste
eller
någon
sådant
med
henne
,
vart
hon
fördenskull
av
rätten
fri
sagt
,
vart
vite
80
mr
på
lyst
att
den
henne
därför
förviter
och
intet
kan
övertygat

Dessa
effterne
är
för
några
år
sedan
komna
till
Ödesheman
,
och
ligger
en
del
av
Åkern
ännu
igen
,
och
felar
efter
utsäde
.

Lasse
Olofsson
i
Aal
tillstod
sig
ha
uppburit
av
h
.
Karins
förre
man
S
.
Olof
skrivare
4
daler
(
på
)
Hökeby
.

Blev
ännu
som
tillförne
dömt
är
Erich
Larssons
barn
i
Mörkarsbo
till
att
njuta
och
behålla
för:ne
Mirkarsbo
för
60
mr
Penningar
både
Jord
och
hus
och
ifrån
Andes
Larssös
barn
som
satt
till
förne
på
samma
hemman
[
Erich
Larsson
i
Fåneby
kärade
till
sin
granne
Pedher
Jönsson
att
han
med
vredesmod
hade
gått
hem
till
honom
och
huggit
honom
i
handen
att
han
där
av
har
evärdligt
Lyte
vart
sack
20
mr
till
treskiftes
och
Målsäganden
12
mr
för
Ljtfhet
,
Item
hade
han
och
slagit
honom
en
blåma
vart
sack
3
mr
och
för
Edsöret
på
hans
Ma:ttz
Nådige
behag
40
daler
.

Men
alldenstund
Michil
Morthesson
bortbytte
3
öres
Land
Jord
mera
än
han
i
Mörkarsboda
bekom
igen
,
skulle
Andreas
Erichsson
som
nu
på
Kätzlinge
bor
betala
Michil
Morthenssons
barn
,
såsom
och
Olof
Matsson
och
hans
Syster
dotter
samma
3
öres
Land
,
efter
som
var
kan
ha
till
att
fordra
.

Så
Allden
Stund
detta
Nu
så
Länge
har
oklandrat
som
be:t
är
,
och
där
Inga
Skäl
och
bevis
hade
där
Något
Att
Fordra
,
Blev
Därför
avsagt
att
be:te
Hans
Humble
skulle
bli
Vid
hemmanet
Efter
Som
tillförne
avsagt
är
,
Och
be:te
Anderss
Matson
och
Jacob
Jnth
:
har
mer
Där
på
tala
som
så
Länge
har
okvalt
Stått
.

Olof
Benchtsson
Benchtz
Son
i
Romstarebo
hade
belägrat
en
knekt
Änka
och
rått
henne
med
barn
vart
sack
3
mr
vilken
är
död
bliven
i
barnsäng
den
där
bekände
för
Ärliga
dannekvinnor
som
då
tillstädes
vore
som
är
h
.
Brita
och
h
.
Kristin
i
Aal
,
att
Olof
var
föga
vållande
där
till
utan
hon
själv
(
hade
lockat
honom
där
till
och
själv
var
orsak
till
sin
död
)
.

Hederlig
och
välLärd
h
.
Andreas
Erici
Kyrkoherde
i
Wendel
Socken
lät
annat
sin
uppbjuda
Holfwebo
hemmanet
det
han
köpt
hade
av
Erich
Joensson
i
Holfwebo
.

Anders
Olofsson
i
Walla
hade
legat
i
Lönskaläge
med
en
knekt
(
sic
)
Änka
h
.
Brita
,
vart
därför
sack
3
mr
.

Kap:
Konungs
Balken
att
böta
Penningar
-
40
mr
för
det
han
smälek
har
talat
om
välborne
Landshövdingen
,
Nämligen
föregivit
att
Anders
Andersson
skulle
ha
givit
Hans
Herlig:t
en
Björnhud
för
det
han
skulle
få
Nämna
till
knektar
Vilka
honom
bäst
Tycktes
,
Vilket
han
och
icke
Neka
kunde
,
Utan
bekände
sig
ha
sådant
sagt
Utav
dåraktighet
,
Uti
sin
stora
fylla
och
druckenskap
.

Noch
avsades
att
Erich
Larsson
i
fåneby
skall
tillställa
Jöns
Larsson
i
Akerby
Uti
Löfstadh
en
halv
spann
Råg
till
,
Uppå
det
Stoköpet
de
sig
emellan
gjort
hade
,
och
ännu
Resterade
.

Såsom
och
fyra
Lass
Äng
Uti
Diupmyran
till
en
behaglig
tid
,
där
om
de
vore
vänligen
förlikta
och
gjorde
varandra
handsträckning
,
att
så
oryggligen
av
dem
båda
hållas
skulle
.

Berättade
och
Befallningsmannen
att
för:ne
Jöns
hade
klagat
på
Jahan
Trostigh
som
fläsket
anammade
,
att
han
skall
ha
vägt
det
bort
,
det
han
icke
eller
bevisa
kunde
,
vart
Jöns
tillsagt
att
betala
fönne
3
få
Fläsk
och
medan
han
och
hade
vitt
andra
där
före
vart
Jöns
sack
40
mr
.

Vart
sagt
att
Matz
skulle
giva
henne
4
'
/
i
daler
gott
mynt
,
och
h
.
Christin
skulle
låta
honom
bekomma
sina
skedar
igen
.

HögLärd
Doktor
Laurentius
Wallius
Tillsporde
rätten
genom
sin
skrivelse
om
han
icke
må
sälja
Erich
Anundsson
det
hemman
i
Granby
som
han
köpt
hade
av
Änkan
h
.
Mariet
som
Lagligen
å
Tingen
år
1630
den
4
November
,
förste
sin
,
år
1631
den
21
Januari
annat
sin
och
samma
år
den
4
Juli
tredje
sin
uppbjudet
och
Lagståndet
är
,
och
tillbjöd
Hans
Vyrdighet
fönne
h
.
Mariet
och
hennes
arvingar
ännu
lossat
och
medan
ingen
var
i
släkten
som
det
lossa
ville
därför
tillsades
Hans
Vyrdighet
Doktorn
att
sälja
vem
honom
täcktes
Äleborna
kärade
till
Akerby
karlarna
att
de
hade
skjutit
ut
vrak
som
drev
in
på
deras
Ängar
,
vart
sagt
att
Akerby
karlarna
skola
En
dag
var
Arbeta
där
på
och
rensa
och
räfsa
samma
vret
tillsammans
igen
,
och
göra
Ängen
rena
vider
bott
där
oftare
klagas
.

Vart
sagt
att
Anders
Höök
och
hans
medarvingar
skulle
behålla
så
länge
den
byggning
räcker
som
han
S
.
fäder
har
där
bygga
låtit
och
icke
längre
,
dock
de
emellertid
där
med
rättvisligen
handla
.

(
1638
)
Den
23
Januari
stod
Lag
ting
i
Wendele
Sockenstuga
uti
Befallningsmannens
Ärlig
och
välbetrodd
Olof
Joenssons
närvaro
dessa
Edsvurna
såtar
i
Nämnden
.

Lars
Morthensson
i
Swartbeckien
vilken
år
1637
den
8
November
fäste
Lag
att
själv
tolfte
göra
sig
fri
för
den
häst
och
föll
som
för
Landsmannen
välaktat
Anders
Högk
är
till
döds
huggna
kom
nu
fram
och
sade
sig
inga
gärningsmän
kunna
bekomma
nu
än
tillförne
,
då
sade
wälb:te
Anders
Hööck
att
där
han
tingat
allenast
en
av
de
Ärliga
män
som
Synade
hästen
,
ville
svärja
med
honom
,
ville
han
där
med
väl
giva
sig
till
frids
,
och
han
skulle
där
med
vara
fri
.

Om
gud
aktig
låter
världen
något
länge
stå
.
så
skola
efter
kommanderne
ingalunda
....
tillåta
....
någon
kvarn
mera
vid
Åbygeby
byggas
.
så
framt
....
ha
sina
ägor
för
skada
behållna
.

Erich
lämnade
detta
till
rättens
omprövande
och
begärde
resolution
här
över
,
med
påstående
,
efter
sin
på
Olof
Olssön
uttagna
stämning
,
det
måtte
han
bli
efter
lag
och
process
bli
ansedd
för
de
håniska
och
skymfliga
ord
,
som
han
utgöt
emot
honom
vid
sista
ting
under
aktionen
med
honom
,
och
pretenderade
expenser
av
Olof
till
24
daler
kopparmynt
för
bägge
tingen
.

timber
eller
gärdsle
;
Ty
hemställs
till
högvälborne
herr
baron
och
landshövdingar
höggunstiga
omprövande
och
förordnande
,
huruvida
vederbörande
må
få
av
allmänningen
hämta
och
hugga
meranämnde
timber
och
gärdsel
med
stör
,
kunnandes
granstockar
brukas
till
stället
och
fourierbostället
väl
behjälpa
sig
,
om
det
får
hälften
av
gärdslet
och
stören
.

Emellertid
tog
sig
rätten
före
att
avhöra
,
vad
dessa
parter
vid
de
övriga
stämningspunkterna
kunna
ha
att
påminna
och
anföra
,
såsom
1:0
vad
soldathusen
angår
,
för
vilkas
behörige
byggnad
Michel
Andersson
erkände
sig
böra
proportionaliter
svara
för
sin
tid
vid
hemmanet
;
även
så
tillstod
han
2:do
sig
vara
på
fördelsspannmålen
skyldig
för
år
1734
2
tunnor
och
för
nästlidet
år
4
tunnor
,
men
att
visa
,
det
allt
vad
av
hemmanet
utgöras
bör
,
/
är
betalat
,
menade
han
vara
tid
nog
till
,
när
vederbörande
låta
förmärka
,
att
de
intet
fått
det
som
av
honom
bör
presteras
.

Beträffande
gärdsgården
så
sade
/
han
,
att
den
var
borta
,
när
han
kom
till
hemmanet
,
änskönt
Lars
Jansson
i
Norrby
intygade
,
att
den
stod
kvar
,
dock
nog
förfallen
,
när
han
år
1720
tjänade
för
dräng
på
Norrby
,
och
att
den
jämväl
var
kvarstående
4
år
därefter
.

Charta
sigillata
penningarna
var
6
daler
24
.
/
.
silvermynt
,
som
vid
detta
ting
i
lådan
influtit
Actum
ut
supra
;
På
tingsrättens
vägnar
A
.
Valtinsson
/
SAKÖRES
LÄNGD
Kronans
Frälsets
Häradets
Målsägandens
Rättens
Drängen
Jonas
Mårtensson
i
Romstarbo
och
kvinnopersonen
Karin
OlofsdoWer
från
Tiärpz
prästgård
böta
för
med
varannan
begått
lönskaläge
,
medan
de
tjänade
tillsammans
på
Hofs
frälsehemman
här
i
socknen
för
två
år
sedan
,
han
10
och
hon
5
daler
silvermynt
samt
stå
sedan
var
för
sig
en
söndags
uppenbara
kyrkoplikt
,
innan
de
absolveras
.
5
5
5
Johan
Ersson
i
Åhrsbo
,
Lars
Mattsson
och
Erich
Andersson
i
Umbärga
,
Michel
Pärsson
i
Myren
,
Lars
Jansson
och
Erich
Ersson
i
Norrby
,
instämde
av
landägaren
Öhrling
,
böta
för
försummat
drevskall
nästWne
5:te
dag
jul
var
sina
6
marker
silvermynt
3
3
3
Michel
Andersson
i
StorEnen
böter
för
3:ne
gånger
försummad
hållskjuts
var
"
sina
3
gånger
3
marker
silvermynt
,
instämd
av
gästgivaren
Ohsengius
i
Läby
.
24
M
Drängen
Erich
Gabrielson
i
Miöhlänge
,
instämd
av
länsmannen
Gabriel
Wretberg
,
böter
,
för
det
han
varit
drucken
,
sina
5
daler
silvermynt
eller
sitter
,
i
brist
av
bot
,
en
söndag
i
stocken
vid
Wändels
kyrka
.
/
2
16
2
16
Bertill
Ersson
i
Massbo
och
soldaten
Erich
Lindberg
böta
,
såsom
contumaciter
uteblir
'
uti
saken
med
hustru
Malin
Berelia
i
Bergby
,
var
sina
2
daler
silvermynt
4
Nils
Andersson
i
Fånby
böter
för
ett
på
Anders
Andersson
ibidem
utgjutit
skälls
ord
sina
3
marker
silvermynt
8
8
8
Summa
4
5
9
11
16
4
2
16
1
Avskrivet
till
till
Kunglige
Hovrätten
.

Det
har
vi
undertecknade
ett
byte
oss
emellan
fastställt
och
gjort
med
de
hemman
vi
här
i
socknen
inneha
,
på
det
sätt
att
jag
,
Pehr
Leufstedt
,
avstår
till
kyrkoherden
här
i
Wändel
,
herr
magister
Erich
Boije
,
mitt
hela
skatte
hemman
i
Gryttby
,
vilket
är
augment
till
rustningsstammen
i
Åkra
,
med
jord
,
hus
och
allt
annat
,
som
därtill
hör
,
tillika
med
Dägare
utjorden
,
Ruddun
dito
med
mera
,
såsom
jag
det
nyttjat
och
innehaft
.

§
.
/
.
kopparmynt
,
dem
min
svåger
Pehr
Niellsson
kvitterat
sig
ha
emottagit
,
återstår
allenast
,
sedan
de
33
daler
kopparmynt
till
den
dels
utlösande
,
som
min
syster
och
Pehr
Niellssons
hustru
Elin
Jansdotter
äger
i
Hökeby
,
bli
avräknade
,
och
den
i:nax
tunnan
råg
antingen
in
natura
eller
med
penningar
blir
betalat
,
femtiotre
daler
kopparmynt
,
varutav
jag
,
Pehr
Niellsson
,
utfäster
mig
att
halvparten
betala
nästkommande
höst
och
den
andra
hälften
hösten
1737
.
/
Som
attesteras
av
Huseby
dnn
2
maj
1736
.

Samma
vret
är
omkring
430
steg
och
nu
är
inlagd
i
gärde
.

Hustru
Eva
tillstod
,
att
hon
slog
bemä
/
de
Nils
Pärsson
med
en
eldtång
över
axlarna
,
för
det
han
var
alltför
otidig
emot
henne
,
med
skällsords
utgjutande
på
henne
av
hora
och
annat
,
samt
beskyllde
henne
för
att
vara
drucken
,
det
hon
dock
likväl
intet
skall
varit
,
men
skall
likväl
intet
tillfogat
honom
någon
åkomma
.

Länsmannen
beropade
sig
alltså
till
vittne
på
drängen
Lars
Ersson
på
Bergby
,
vilken
till
vidare
utan
ed
berättade
,
det
Nils
Pärsson
,
som
låg
hos
honom
i
sängen
,
skall
först
kallat
dottern
i
gården
FyllCatrina
,
och
när
hustru
Eva
därpå
svarade
,
alla
kallar
Ni
fulla
,
skall
han
även
många
gånger
kallat
henne
FyllEva
.
/
Sedan
de
således
länge
hade
kivat
med
skällsords
utgjutande
på
var
annan
och
Nils
Pärsson
sagt
,
att
hon
var
en
hora
samt
att
soldaten
Lindberg
var
hennes
horekamp
,
skall
Eva
sport
honom
till
,
om
han
det
tillstå
kunde
,
och
emedan
han
än
då
intet
vände
igen
med
skällsord
på
henne
,
skall
hon
tagit
till
en
eldtång
och
slagit
honom
med
,
där
han
låg
i
sängen
,
några
slängar
,
varför
han
skall
sprungit
opp
utur
sängen
till
matmodern
och
bett
henne
se
,
hur
hustru
Eva
hade
slagit
honom
,
var
på
han
skall
föst
henne
utur
stugan
och
gjort
ett
fasligt
alarm
,
vilket
skall
föranlåtit
Lars
Ersson
till
att
gå
opp
utur
sin
nattsäng
och
fråga
dem
till
,
vad
de
hålla
för
ett
väsende
,
samt
bedja
Nils
betänka
,
vad
han
gjorde
,
och
gå
till
sängs
igen
.

Olof
Olssön
beropade
sig
likafullt
på
sin
och
sina
förfäders
gamla
hävd
och
de
vid
första
tinget
härom
producerade
attester
,
den
han
förmenade
sig
böra
få
till
godo
njuta
,
till
dess
han
blir
lagligen
dömd
ifrån
bemä
/
de
hävd
och
vägs
nyttjande
;
varandes
nöjd
med
att
i
mellertid
få
köra
över
ängen
,
dock
intet
vidare
än
när
han
någon
gång
kan
ha
nödigt
att
fara
där
över
till
allmänningen
och
Tiärpz
kvarnar
med
sin
mäld
,
vilket
,
såsom
ovanförmält
är
,
protesterades
av
svaranden
,
med
sin
expensräknings
insinuerande
på
81
daler
8
.
/
.
kopparmynt
för
alla
tingen
.

Och
vad
ärtesåningen
angår
,
så
skall
den
skett
därav
,
att
Brundin
på
Ohsengii
begäran
,
emot
det
att
han
skulle
participera
med
honom
uti
extraordinarie
utgifterna
,
stängt
in
ett
stycke
åker
åt
honom
till
att
med
ärter
beså
,
men
emedan
det
intet
skedde
,
skall
han
besått
bemälde
åkerstycke
med
ärter
och
själv
betalat
extraordinarie
utgifterna
.
5:to
ville
han
ha
ersättning
av
Ohsengiws
,
för
det
han
skall
tagit
tvenne
åkerstycken
av
hemmanet
och
givit
åt
en
torpare
;
skolandes
han
6:to
intet
tagit
emot
något
rov
eller
ärtelands
gärdsel
,
när
han
kom
till
hemmanet
,
mindre
fört
något
därifrån
,
utan
stängt
opp
det
han
huggit
på
Grytby
skog
,
där
det
behövts
vid
hemmanet
.

Å
ryttmästarens
välborne
herr
Thomas
Rudebecks
vägnar
anhöll
kyrkoherden
ärevyrdige
och
höglärde
herr
magister
/
Erich
Boije
om
denna
rätts
attestatum
,
hur
vi
då
bemälde
herr
ryttmästares
eller
dess
kära
husfrus
frälsehemman
,
fyra
i
Karby
och
ett
i
Åhsbo
här
i
soclnen
belägna
,
är
med
någon
inteckning
eller
på
något
annat
sätt
här
vid
rätten
graverade
,
var
på
till
efterrättelse
och
behörig
säkerhet
lämnades
,
det
bemälde
hemman
är
varken
med
någon
inteckning
eller
på
något
annat
sätt
här
vid
rätten
besvärade
utan
alldeles
fria
och
lediga
därifrån
.

Responsum
,
8
dagar
,
samt
att
han
,
medan
sjukdomen
påstod
,
intet
låg
stadigt
utan
låg
ibland
till
sängs
,
ibland
gick
han
oppe
,
skolandes
ännu
intet
vara
bättre
fri
därifrån
,
än
att
han
alltsomoftast
har
brytningar
av
samma
sjukdom
,
varförutan
han
också
skall
vara
så
svag
till
sitt
huvud
,
att
han
ibland
raglar
på
sned
,
utan
att
han
just
är
sjuk
.

Erich
Andersson
,
att
Ekeroth
den
tiden
uti
nästlidna
fasta
,
när
snön
begynte
gå
bort
,
var
hos
honom
till
att
sömma
skor
men
skall
av
frossan
så
blivit
betagen
,
att
han
intet
förmåde
göra
något
arbete
utan
nödgades
gå
hem
,
vilket
skall
kontinuerat
med
honom
hela
våren
,
jämte
bröstsjuka
.

Quasstio
till
Ekeroth
,
vi
han
intet
höll
sig
från
bränn
vin
emellan
predikningarna
,
när
han
visste
,
att
han
var
så
svag
till
att
det
kunna
tåla
?

Sammaledes
presenterades
och
upplästes
det
bytes
brev
av
den
19
juli
innevarande
år
,
som
välborne
herr
Carl
De
Geer
igenom
inspektorn
herr
Erich
Touschier
slutit
och
fastställt
emellan
sig
och
nämdemannen
Anders
Andersson
i
Libbarbo
och
dess
son
Bängdt
/
Andersson
,
av
dem
underskrivet
samt
till
vittnes
av
inspektorn
herr
Gustaf
Kiörning
,
varmedelst
välbemälde
herre
till
honom
,
Anders
Andersson
,
uppdraget
skatträttigheten
av
det
hemman
i
Walla
,
som
sonen
Bengt
Andersson
hit
tills
brukat
såsom
dess
frälses
landbo
,
och
under
samma
hemman
jämväl
få
äga
och
nyttja
utjordarna
,
Wibbelbohle
och
Wallaboda
kallade
,
den
förra
om
sex
och
den
senare
om
tolv
penningland
,
varemot
Anders
Andersson
avstått
sitt
skatte
hemman
,
Stor-En
kallad
,
även
här
socken
beläget
,
bestående
av
4
.
/
.
land
med
allt
vad
som
där
till
hör
,
såsom
det
nu
befinns
och
för
ögonen
står
,
samt
där
till
av
ålder
lytt
och
legat
har
,
tillägnandes
detsamma
herr
Carl
De
Geer
att
därmed
disponera
och
råda
som
all
annan
sin
lag-
och
välfångade
egendom
;
I
följe
varav
blev
,
uppå
notarien
Hoffmans
anhållan
,
bemälde
StorEns
hemman
,
med
alla
/
dess
tillhörigheter
,
välborne
herr
Carl
De
Geer
tillhanda
uppbjudit
första
gången
.

Denna
skuld
erkände
Anders
Jansson
till
48
daler
kopparmynt
,
det
övriga
disputerade
han
såsom
efter
dess
mening
för
mycket
honom
påfört
för
en
häst
,
den
han
sade
sig
ha
av
inspektorn
Hagel
bekommit
;
men
sedan
han
blev
av
dess
bok
underrättad
om
skuldens
riktighet
,
så
kunde
han
den
intet
frångå
,
varför
och
emedan
befallningsmannen
välbetrodde
Philip
Befwert
lovade
sig
så
skola
laga
,
att
den
skall
vid
Tobo
efter
hand
bli
betalat
,
och
inspektorn
Hagells
fullmäktig
,
sonen
gruvfogden
Carl
Hagel
,
var
där
med
nöjd
,
allenast
han
också
får
ovannämnde
expenser
av
honom
;
/
Alltså
förblir
det
ock
där
vid
,
dock
så
,
att
Anders
Jansson
jämväl
bör
uti
expenser
till
inspektorn
Hagel
erlägga
6
daler
kopparmynt
.

Inspektorn
herr
Erich
Hagell
hade
också
instämt
följande
för
skuld
till
sig
,
nämligen
Jan
Andersson
i
Hålfwarbo
,
nu
i
Botarbo
,
om
90
daler
,
Jan
Pärsson
i
Råssla
om
84
daler
och
Erich
Olssön
i
Myrstugan
eller
Fånby
om
71
daler
5
.
/
.
kopparmynt
,
dem
han
fördenskull
av
dem
ville
ha
,
med
expenser
till
14
daler
8
.
/
.
kopparmynt
av
dem
vardera
,
betalade
.

Och
som
hygget
,
efter
bemälde
rors
anledning
,
där
inom
skall
vara
skett
,
så
förmenade
han
,
det
de
böra
lämnas
otilltalade
därför
.

Klagades
ock
mycket
av
hela
församlingen
,
men
besynnerligen
av
frälse
Inspektorn
J
.
C
.
Kralle
över
det
stora
oljud
och
oväsende
,
som
*
se
Inledning
.
!
)
se
Noter
.

Flickan
tillspordes
:
om
hon
all
ovan
anförda
tjuvnad
begått
hade
?
varpå
hon
svarade
:

Hon
visste
ock
icke
det
ringaste
för
sin
odygd
skämmas
:
mindre
om
förlåtelse
bedja
,
utan
med
fräcka
gebörder
skickade
och
tedde
hon
sig
för
allas
ögon
.
§
8
.

Angav
Eric
Larsson
uti
Låskebohl
,
hur
mjölnarhustrun
uti
Wallbyqwarn
,
utan
rättighet
alltid
tränger
sig
in
,
uti
dess
Hustrus
och
Bänkkamrats
Stolrum
i
kyrkian
,
och
icke
allenast
dem
tränger
,
utan
ock
föregav
,
att
de
till
bänkrummet
berättigade
ofta
uteslutna
bli
.

Antyddes
ock
Församlingen
,
hur
General
Löjtnanten
,
högvälborna
Herr
Baron
Eric
Fitinghoff
begär
och
påstår
:
det
måtte
Nedergården
uti
Biurstorp
hädanefter
höra
till
Biurstorpa
Roote
och
icke
till
Båltznääs
Roota
;
emedan
på
den
tiden
,
då
åtskilliga
ägare
varit
till
Juhla
och
Dufweholms
Säterier
,
är
gårdarna
uti
Biurstorp
,
och
blev
delade
till
åtskilliga
Rootar
;
vilket
ock
alla
fann
för
skäligt
att
stadsfästa
.
§
3
.

Påmindes
och
angavs
hur
Skräptorpa
Gossar
,
tillika
med
gossen
ifrån
Sömmerskestufwan
,
gjorde
oljud
på
Bönedagen
och
övade
Stim
på
Kyrkovallen
under
Högmässo
Gudstjänsten
.

Så
vara
slutat
och
avgjort
,
attestera
,
Anno
die
et
loco
,
ut
supra
.

Närvarande
barnets
morbroder
i
Tyble
,
Nils
Nilsson
i
Tyble
,
utfäste
å
sin
faders
vägnar
,
att
barnet
hos
sin
morfader
skulle
njuta
sin
uppfostring
,
och
blev
så
därpå
enhälleligen
beviljat
,
att
barnet
undfå
skulle
faderns
fattigdel
,
som
ett
allmosehjon
utom
fattighuset
,
men
icke
där
intagas
.
§
10
.

Item
tillspordes
:
om
Församlingen
än
vidare
förskott
göra
ville
efter
den
förra
antagna
metoden
,
att
nämligen
)
av
var
person
,
som
begick
Herrens
Heliga
Nattvard
,
ung
eller
gammal
,
skattlagd
eller
oskattlagd
)
skulle
årligen
erlägga
16
.
/
.
kmt
,
tills
Klockan
blev
betalad
:

Häruppå
gav
de
närvarande
herrskapen
,
med
betjänter
och
menige
man
,
sina
otvungna
vota
till
Ryttaren
Anders
Jenzell
,
såsom
den
tjänligaste
och
skickligaste
.
5
2
.

Ropades
fram
man
ifrån
man
,
och
by
efter
by
i
församlingen
/
:
för
de
bortavarande
svarades
och
gjordes
redo
av
Roota
mästarna
och
Sexmännen
:
/
att
efter
Maxime
)
Venerandi
)
Consistorii
)
av
d
.
25
febr
:

Sistlidne
)
utgångna
skriftliga
befallning
,
det
skulle
ifrån
alla
församlingar
berättelse
tidigt
inflyta
,
hur
många
barn
lärt
läsa
i
bok
,
eller
därmed
börjat
och
begynnt
ifrån
Riksdagen
1723
till
1727
,
och
ifrån
1727
till
innevarande
år
;
var
och
en
för
sig
och
sina
barn
,
skulle
sig
härom
utlåta
och
redogöra
.

Skärptes
vederbörligen
)
den
vederstyggliga
osed
och
vanart
,
som
somliga
uppenbarligen
bevisa
,
med
sitt
otidiga
)
tobaksrökande
uti
KlockarKammaren
,
besynnerligen
före
allmänna
Gudstjänsten
och
innan
Sammanringningen
;
och
som
detta
tillförende
en
gång
blivit
föreställt
,
men
ingen
verkan
haft
,
uppläste
Pastor
Kungl.
Förordningen
de
anno
1714
d
.
25
Martii
,
som
vid
böter
förbjuder
att
röka
tobak
vid
kyrkorna
på
Helgdagarna
.

Några
som
suttit
uti
Socknens
Gravkapell
sade
sig
väl
det
samma
hört
,
då
de
efter
klockslagen
hört
eller
tyckt
,
att
någon
av
de
vanartiga
barnen
på
backen
måtte
ha
hanterat
klocksträngen
,
ville
ock
ha
gossen
i
Sömmerskestugan
suspekt
)
Men
ehuru
Pastor
förmanade
,
att
man
skulle
detta
uttryckligen
uppenbara
,
fanns
dock
ingen
,
som
tillförlitlig
underrättelse
härom
giva
kunde
.
§
6
.

Item
Resol
.
på
allmogens
besvär
1720
§
41
uppläst
var
,
av
innehåll
att
oskattlagda
Torpare
så
väl
som
inhyses
hjon
,
även
de
som
sitta
i
Backstugor
,
skola
i
Prästegårds
Byggnad
participera
:
påstod
församlingen
enhälligt
,
att
likmätigt
denne
Kungl.
Förordningen
,
ovannämnde
Församlingens
invånare
,
skulle
till
Byggnaden
proportionaliter
biträda
.
§
9
.

Framkallades
tjänstegossarna
ifrån
Stenstorp
,
Gatubohl
och
Olofstorp
,
som
emot
förra
träffade
beslut
,
hade
förmaningar
att
sitta
bak
i
kyrkan
och
på
läktaren
att
göra
förargelse
,
buller
och
stim
;
och
dömdes
tjänstegossarna
ifrån
Stenstorp
,
att
sitta
nästa
söndag
i
Stocken
,
men
de
andra
gossarna
befriades
ifrån
straffet
denna
resan
,
med
allvarsam
förmaning
.
§
10
.

Men
alldenstund
församlingens
ledamöter
själva
veta
att
en
del
av
dem
är
tröga
och
tredska
,
i
rättan
tid
ifrån
sig
avgiva
det
som
på
Sockenstämmorna
till
kyrkans
reparation
och
andra
förnödenheter
frivilligt
slutet
blivit
,
så
begärdes
och
påstods
av
de
närvarande
enhälligt
,
att
i
den
händelse
icke
alla
villigt
och
enhälligt
,
med
betalningen
sig
inställde
på
förbemälta
tid
,
måtte
man
höga
landshövdinga
ämbetet
i
ödmjukhet
anlita
,
om
nådig
handräckning
:
på
det
att
det
åbelöpande
Intresset
varken
måtte
flera
år
erläggas
,
icke
eller
de
villiga
att
betala
,
med
mera
onödig
utgift
,
för
de
tröga
och
tergiverserandes
skuld
,
graveras
)
§
3
.

Men
emedan
besynnerlig
2ne
var
,
som
i
de
förra
åren
alltid
tredskat
,
dem
Kyrkoherden
för
denna
gång
ej
heller
ville
utnämna
,
ty
blev
de
ock
förmanade
till
bättre
besinnande
av
ett
så
angeläget
verk
.

Församlingen
tog
denna
sak
uti
vederbörligt
betänkande
,
och
alldenstund
församlingens
samtliga
Respektive
Herrskap
,
skriftligen
sitt
goda
jaord
där
till
på
Sockenstämman
ingivit
,
blev
slutet
endräktligen
,
att
samma
lille
inkomst
av
församlingens
fria
villa
,
Komministern
årligen
tillflytta
skall
uti
dess
tjänstetid
,
dock
utan
att
detta
efter
honom
,
dragas
må
till
en
vana
,
eller
Församlingens
tunga
.
§
17
.

Likaledes
påstod
Sexmannen
för
Måsstorpa
Roota
,
Pär
Andersson
i
Remmerööstorp
,
orlof
och
blev
så
efter
honom
till
Sexman
kallad
unga
Lars
i
Biörnkällan
,
men
skulle
han
,
såsom
då
frånvarande
,
samma
syssla
ej
vilja
sig
åtaga
,
föll
man
på
Lars
Pehrsson
i
Kåhlberga
,
som
då
tillstädes
var
.

Härtill
kunde
man
icke
samtycka
,
i
någondera
måtto
,
förr
än
Gabriel
kunde
skaffa
sig
fulla
bevis
till
sin
talan
,
då
man
sedermera
ville
giva
ett
visst
svar
,
hänvisande
man
Gabriel
till
laga
Forum
,
om
han
förmenar
sig
vara
av
Claes
uti
sin
tillständiga
Rätt
förfördelat
.

Framträdde
förlovade
soldaten
Lars
Stenbom
,
och
uti
sin
stora
nöd
och
brist
,
begärande
av
församlingen
någon
assistans
av
de
fattigas
Kassamedel
,
att
betala
de
medikamenter
med
vilka
Stadsfältskären
uti
Nycköping
Herr
Wilhelm
Zachrisson
,
förmedelst
Guds
Välsignelse
hjälpt
honom
ifrån
sin
svåra
Gangrena
och
värk
i
dess
högra
hand
,
emedan
han
själv
ej
hade
något
där
till
att
använda
.

Som
Assessorskan
Välborna
Fru
Florentina
Hildebrand
på
Erichsberg
,
har
av
den
6
juli
sistlidne
skriftligen
vid
handen
givit
,
det
hon
fordrar
dagsverken
av
Oxlegården
och
Sömmerskestugan
,
vilka
små
lägenheter
härtills
varit
Komministern
uti
församlingen
,
ärevördige
och
Vällärde
Herr
Georg
Netzelius
till
disposition
anslagen
av
salig
)
framlidne
Greven
och
lagmannen
Herr
Carl
Adolph
Gyllenstierna
alldenstund
dessa
lägenheter
är
fru
Assessorskan
,
uti
dess
Jordebok
,
utan
något
förbehåll
,
under
sådan
titel
uppförde
:

Men
förbehöll
sig
församlingen
att
icke
framledes
graveras
med
denna
fattigstugas
vidmakthållande
,
emedan
den
ordinarie
socknens
fattigstuga
,
för
dess
räkning
och
ansvar
står
;
Varpå
bifölls
,
att
denna
lilla
Stugan
alltid
bör
med
fattigkassans
propra
medel
,
under
och
vidmakthållas
.

Utlovade
Församlingen
,
att
strax
efter
Andetiden
,
med
spanande
förfärdiga
den
andelen
av
norra
Kyrkotaket
,
som
ännu
ofärdigt
är
.
§
8
.

Föreställdes
i
sammankomsten
,
Eric
Siggesson
i
Ramsiöhult
,
som
förfallolös
på
4
års
tid
uteblivit
ifrån
de
ordinarie
Catechismi
förhören
samt
sista
åren
icke
eller
tillhållit
sina
2
söner
att
sig
infinna
;
Påståendes
Kyrkoherden
,
att
han
efter
Kungl.
Kyrkolagens
2
Gap
:
och
9
§
m
)
skulle
plikta
till
kyrkan
28
.
/
.
smt
.
men
som
bemälte
Eric
Siggesson
gjorde
offentlig
avbön
,
,
samt
gjorde
försäkran
om
verklig
ändring
,
blev
honom
plikten
,
under
allvarsam
förmaning
,
denna
resan
tillgiven
.
§
6
.

Lovade
ock
församlingen
,
att
nästkommande
Söndag
,
vill
Gud
,
giva
ett
ändligt
svar
,
om
det
sätt
och
expedient
på
vilket
den
vansinniga
änkan
uti
Nordanås
skall
uti
församlingen
bli
underhållen
,
emedan
man
icke
kan
henne
uti
sockenfattigstugan
vårda
.
(
Se
vidare
prot
.
28
/
10
1734
,
§
4
)
.

Kontinuerades
med
den
påbegynta
Stolläggningen
,
så
uti
HuvudKyrkan
som
GravKapellet
,
både
med
de
ordinarie
så
väl
som
de
kallade
Rootstolarna
,
och
kom
man
därmed
uti
enighet
och
gott
överenskommande
,
till
ett
ändligt
slut
,
som
StoldelningsInstrumentet
utvisar
.
§
2
.

Så
ock
att
den
gamla
)
och
sjukliga
Olof
i
Hälletorp
,
måtte
av
församlingens
fattigas
andel
,
uti
kost
och
penningar
,
njuta
så
stor
del
,
utom
fattigstugan
,
som
den
avlidne
Jöns
Sarfwe
i
Nästorp
,
förr
njutit
.

Anno
1735
den
1
Maj
,
blev
på
Alman
Valborgsmässo
SockenStämma
,
följande
avslutat
.
$
1
.

Avslutades
,
att
Eric
Larsson
ifrån
Låskebohl
,
Bengt
Persson
ifrån
Kåhlberga
,
Per
Månsson
ifrån
Sundstufwan
,
Anders
Thomsson
ifrån
Råstock
,
hädanefter
skola
del
njuta
av
de
fattigas
förskott
,
utom
fattighuset
,
så
ock
den
gamle
)
Michel
ifrån
Kåppartorp
,
som
fick
tillstånd
att
ha
husrum
uti
nya
fattighuset
,
med
den
del
av
underhåll
,
han
tillförende
njutit
,
men
icke
mera
för
denna
gången
.

Utlovade
Församlingen
,
att
innan
andetiden
infaller
,
med
spanande
förfärdiga
den
andelen
av
norra
Kyrkotaket
,
som
ofärdig
är
;
vartill
för
Kyrkans
medel
är
köpt
Spån
,
och
av
Erstorpa
och
Dahls
Rootar
,
nederkört
till
Kyrkan
ifrån
Fäboda
,
för
3
dagsverken
räknat
vart
lass
.
§
7
.

Kom
Församlingens
invånare
därom
överens
,
att
uti
instundande
Vinter
betala
till
Kyrkan
igen
de
penningar
och
medel
,
som
Snickaren
och
Smeden
fått
i
betalning
av
Kyrkan
för
Stol
och
BänkArbetet
,
nämligen
2
dr
12
.
/
.
kmt
på
vart
skattlagt
matlag
.

Upplästes
det
förra
och
nästledna
ValborgsmässoSockenstämman
hållna
Protokoll
,
som
till
alla
delar
vidkändes
.
§
2
.

I
övrigt
utfäste
sig
ock
Församlingen
,
att
vid
samma
tillfälle
vilja
erlägga
till
små
spiks
upphandlande
,
på
stollistorna
1
.
/
.
kmt
av
var
Person
,
som
för
sig
betalar
till
Stolrummet
.

Begärandes
att
med
samma
slags
tak
,
på
den
ännu
ofärdiga
ringmuren
skulle
kontinueras
för
mindre
omkostnad
skuld
.

Valdes
till
Kyrkovärd
,
med
enhälligt
omröstande
av
hela
Församlingen
,
Pehr
Pehrsson
uti
Prästorp
,
uti
den
avlidne
Nämndemannen
och
Kyrkovärden
Carl
Bengtssons
ställe
i
Walla
,
dock
med
det
förbehåll
,
att
bemälta
Carl
Bengtssons
änka
,
skulle
pro
anno
1735
,
njuta
och
behålla
dambspann
§
6
.

Joen
förklarade
sig
ha
mycket
illa
gjort
och
utlovade
bättring
.

Tillsades
församlingen
,
att
i
Vinter
framskaffa
brädor
och
Spån
,
som
restera
till
det
påbegynta
Ringmursarbetet
,
emedan
uti
innestundande
Vår
,
om
Gud
vill
,
man
åter
ett
stycke
av
ringmuren
skall
företaga
att
reparera
,
efter
samma
sätt
och
vis
,
som
det
redan
förfärdigade
skett
har
.

Även
berättade
ock
Simon
:
att
vid
påfordran
,
skall
han
för
sig
kunna
utvisa
sagsman
till
sådant
rykte
.

Uppvisade
också
ett
Malmströms
brev
,
därutinnan
han
debiterar
Kyrkoherden
för
mindre
samvetsgrann
,
om
arbetet
ej
bättre
anses
och
betalas
skulle
,
än
som
projekterat
var
uti
Församlingens
sammankomst
,
till
600
daler
kmt
,
och
någon
diskretion
.

§
.
Byggninga
)
Balken
stadgar
om
allmänna
hus
Byggnad
,
och
dagverken
därtill
;
så
att
på
det
arbetet
icke
skulle
bli
för
långsamt
,
om
dagverken
allenast
efter
hemmantalet
göras
skulle
,
de
samma
av
vart
matlag
presteras
borde
,
de
oskattlagda
härifrån
undantagna
;
samt
att
därmed
begynnas
borde
uti
Foglöö
Roota
,
därest
dagverksordning
och
omgångar
sist
stannat
hade
.
§
5
.

Vid
samma
tillfälle
,
ställdes
även
flera
gossar
för
ögonen
deras
slemma
vanart
vid
allmänna
Gudstjänstens
förrättande
,
nämligen
Eric
Jonsson
i
tjänst
vid
Kåhlgölet
,
den
avlidne
Jonas
Wallgrens
son
,
förty
han
hade
suttit
kvar
i
Fattigstugan
,
när
Gudstjänsten
påstod
,
som
Sexmannen
i
Heden
visste
att
berätta
;
Föravskedade
nummersoldaten
Arenberg
son
,
Anders
vid
samma
namn
,
tjänande
hos
Anders
Larsson
i
Remmeröö
,
vilken
Kyrkoherden
funnit
stående
på
Kyrkobacken
,
även
under
påstående
Gudstjänst
,
vid
anresande
Folks
förvägnar
;
Så
ock
gästgivaren
Emanuel
Stålts
Tjänstegosse
uti
Stensiö
Johan
Bengtsson
vid
namn
,
vilken
stått
utan
för
Kyrkodörren
,
och
icke
velat
gå
därin
under
Predikan
.

Uppå
Kyrkoherdens
tillfrågan
:
om
Församlingen
kunde
giva
något
förslag
på
någon
tjänlig
Socken
Skomakare
,
uti
Olof
Larssons
ställe
som
antagit
Krigstjänst
och
bort
marscherat
:
svarades
,
att
de
icke
nu
visste
någon
skicklig
att
föreslå
;
men
Välborne
Herr
Ryttmästare
Hildebrand
behagade
vara
så
god
,
och
lovade
göra
Socknen
den
hjälp
och
Tjänsten
att
försöka
om
icke
möjligt
vara
kunde
,
förmå
någon
av
sina
hantverkare
vid
sina
utom
denna
orten
belägna
Säterier
,
att
flytta
hit
upp
.

Så
beslöt
Församlingen
,
att
av
de
övriga
7
Rootar
,
låta
leverera
50
st.
Tak
Torv
på
vart
helt
hemman
;
befinnandes
sig
invånarna
uti
de
större
Byar
och
gårdar
nedan
vid
Kyrkan
,
villiga
att
ändå
mera
Torv
framskaffa
,
om
behövas
skulle
,
och
vid
annat
tillfälle
njuta
vedergällning
på
dagverken
,
etc.
emot
de
andra
Rootar
,
som
obekvämare
ha
slika
varor
att
framskaffa
,
samt
uti
samma
7
Rootar
att
avgiva
2
st.
Bräder
på
vart
helt
hemman
och
proportionaliter
på
de
mindre
,
vilket
gör
ungefär
9
toffter
och
några
bräder
,
kunnandes
man
de
bräder
som
överskjuta
,
till
ett
annat
behov
och
tarv
förvara
.

Således
vara
avslutat
och
avhandlat
,
Betyga
på
Församlingens
vägnar
J
.
Dalenius
PL
.

Klagade
Per
Persson
uti
Högen
högeligen
däröver
,
att
i
förledne
sommar
skall
honom
på
dess
förfäders
gravplats
skett
orätt
och
förnär
,
då
Kårtorpa
bårlag
därjämte
grävt
,
påståendes
sådant
måtte
bli
behörigen
rättat
;
Kyrkoherden
förmodade
väl
sådant
icke
skett
av
någon
med
uppsåt
och
vilja
,
men
håller
det
förehava
kunna
lätteligen
skett
av
våda
,
emedan
kyrkogården
är
ganska
liten
och
trång
,
förmanade
därför
församlingen
,
att
vid
de
tillfällen
,
som
de
för
sina
döda
gräva
,
all
möjlig
aktsamhet
brukas
måtte
,
att
på
de
nästbelägna
lägerplatser
ingen
skada
ske
måtte
.
§
13
.

Juli
,
inkallades
Församlingen
uti
Sockenstugan
efter
sluten
Gudstjänst
,
då
Plurimum
Venerandi
Consistorii
Cirkulär
skrift
under
d
.
29
Juni
sistfallne
,
kungjordes
,
av
följande
innehåll
;
Konsistorium
vill
ha
kungjort
,
att
emedan
på
domkyrkans
bekostnad
,
Tryckeriet
därsammastädes
,
är
med
kostliga
nya
stilar
försett
,
varpå
man
prov
längesedan
lämnat
,
och
Boktryckaren
Lars
Collin
utlåter
sig
vilja
lägga
upp
Psalmböcker
på
gott
papper
,
allenast
för
1
dr
8
.
/
.
kmt
Exemplaret
;
ty
begäres
att
som
Församlingarnas
respektive
ledamöter
utan
tvivel
behöver
Psalmböcker
för
sig
och
sina
barn
,
det
herrar
Pastores
nu
genast
var
i
sin
församling
ville
uppbära
penningar
,
eller
av
Kyrkans
medel
prenummerera
till
så
många
Exemplar
,
som
åstundas
,
samt
medlen
tillika
med
Specifikationen
därpå
,
igenom
herr
Probsten
,
med
det
första
till
Konsistorium
överstyra
,
kunnandes
man
försäkra
,
att
Exemplaren
inom
ett
års
förlopp
skola
få
av
hämtas
,
då
Psalmboken
kan
has
för
sju
ringare
pris
än
eljest
,
och
kyrkorna
icke
desto
mindre
,
återfå
den
prenumererade
summan
med
därpå
löpande
Intresse
.

Församlingen
stannade
i
det
slutet
:
att
ehuru
väl
många
i
socknen
kunde
under
närvarande
svåra
tider
,
behöva
längre
denna
Krediten
av
Kyrkan
,
dock
likväl
till
att
undvika
den
olägenheten
,
att
enär
vid
hemmanen
ömsas
åboar
,
den
tillträdande
icke
måtte
komma
att
betala
,
vad
den
avträdande
lånat
,
blev
enhälleligen
slutat
,
att
Pastor
till
Sexmännerna
,
en
var
i
sin
Roota
,
skulle
listor
utlämna
,
varefter
dessa
penningar
må
inkasserade
varda
.
§
3
.

Vad
det
angår
,
som
skulle
någon
under
sken
vilja
göra
sig
berättigad
att
rubba
de
i
KyrkoKoret
belägna
och
förmälda
gravarna
,
eller
någon
grift
för
sig
därstädes
reparera
,
så
lär
ej
någon
vara
av
ett
slikt
Sinnelag
;
men
beträffande
det
att
fröken
protesterar
emot
Stolrums
byggande
på
mer
omnämnda
Jula
grifter
,
så
lär
det
så
mycket
mindre
gälla
,
som
ej
allenast
i
denna
Kyrka
,
utan
ock
allestädes
brukligt
är
,
att
på
gravar
bygga
bänkar
och
Stolrum
.
§
12
.

Således
vara
avhandlat
,
betyga
på
Församlingens
vägnar
:

Föreställde
Kyrkoherden
Församlingen
den
slemma
vanart
han
kommit
i
erfarenhet
om
,
att
uti
Fattigstugan
,
skall
nu
åter
börjas
med
brännvinssäljande
på
Sön
och
högtidsdagar
,
emot
de
förr
kungjorda
Kungl.
Förbud
och
förordningar
,
med
mera
,
/
:

Härpå
svarades
:
att
ehuru
hela
Församlingen
hade
sig
förmodligen
bekant
,
det
uti
sådana
Kyrkomål
,
man
alltid
,
så
väl
som
i
alla
andra
tillfällen
,
har
haft
avseende
på
de
fattiga
,
och
denne
avgiften
icke
alltid
till
det
strängaste
av
dem
utfordrat
,
synes
likväl
betänkligt
,
att
alldeles
denna
lilla
avgiften
för
Kyrkan
,
som
är
en
Pupill
och
har
städse
många
oundgängliga
tarvor
,
indraga
,
helst
den
icke
bör
anses
annorlunda
,
än
som
en
skyldig
och
kristlig
erkänsla
mot
Gud
och
Hans
Heliga
Hus
,
den
kyska
Brudar
villigt
borde
erlägga
,
såvida
deras
förmåga
någorlunda
det
tillåter
,
därför
att
Gud
dem
i
alla
deras
livsdagar
bevarat
för
skada
och
skam
på
deras
goda
namn
och
ärliga
rykte
med
mera
:

Klagade
Socken
Skräddaren
Sven
Svensson
över
Jöns
Larsson
i
Björnmogen
att
han
förfördelat
honom
med
syende
uti
Walla
by
,
samt
att
det
samma
skall
honom
ofta
ske
av
Nummer
)
Soldaten
)
Lars
Snack
och
avskedade
Lars
Norman
,
vilka
även
skola
ha
gossar
med
sig
,
när
de
göra
församlingen
tjänst
.

Herr
Löjtnant
Lidstrand
tilltalade
Jöns
Larsson
allvarsamt
,
med
befallning
att
bruka
hemmanet
,
och
låta
bli
Skräddarhantverket
och
angående
de
senare
,
så
är
tillförne
av
Kungl.
Förordningen
kunnigt
,
att
nummersoldater
,
när
de
hemma
vistas
vid
sina
boställen
,
utan
tilltal
äga
frihet
att
idka
sina
hantverk
,
men
icke
ha
tillstånd
att
betjäna
sig
av
lärogossar
;
Vilket
tillsades
Sexmännen
att
göra
dem
å
Församlingens
vägnar
kunnigt
,
alldenstund
de
icke
tillstädes
var
.
§
24
.

Nils
Nilsson
i
Remna
Per
Persson
i
Stensjö
Nämbdeman
kyrkovärd
Anders
Andersson
i
Foglöö
sexman
Anno
1744
den
21
October
,
höll
man
efter
föregången
vanlig
pålysning
,
allmän
Mickelsmässo
SockenStämma
med
St.
Malms
Församling
uti
närvaro
av
respektive
och
Välborne
herrskapet
på
Ericksberg
med
de
övriga
respektive
Församlingens
herrskapers
Betjänter
,
samt
Församlingens
Kyrkovärdar
,
Sexmän
,
äldste
och
menige
man
,
då
följande
blev
föreställt
och
avhandlat
.
§
1
.

Häruppå
projekterade
Kyrkoherden
:
att
om
Församlingen
ville
påtaga
sig
att
Spana
sin
del
av
Taket
,
vartill
ungefärligen
skulle
betarvas
Tio
tusen
spån
å
15
dr
,
gör
150
dr
,
även
så
mycket
spik
å
9
dr=90
dr
kmt
,
sex
Tolfter
Bräder
å
6
dr
gör
36
dr
samt
provisionaliter
till
Byggmästaren
30
dr
eller
40
,
alt
i
Kopparmynt
,
gör
en
Summa
av
318
dr
vid
pass
,
mer
eller
mindre
:

Samma
avgift
påstod
ock
Olof
Larsson
sig
årligen
böra
undfå
av
Anders
Jönsson
uti
Markstugan
;
vilket
Församlingen
prövade
skäligt
,
så
vida
Anders
Jönsson
nu
frånvarande
,
åstundar
obehindrat
samma
hantverk
hädan
som
härtills
idka
.
§
11
.

En
och
annan
i
Församlingen
,
såsom
Simon
Larsson
uti
Afrad
med
flera
,
ville
påstå
,
att
den
så
kallade
Brudstadsgången
skulle
alldeles
upphävas
och
avskaffas
;
Men
målet
blev
;
med
de
flera
,
till
nästa
ValborgsmässoSockenStämman
,
vill
Gud
!
uppskjutet
.

Berättade
även
Kyrkoherden
,
att
han
nödgats
i
Stockholm
förackordera
en
annan
Bleckslagare
,
till
Klocktornets
betäckande
,
än
den
i
förstone
betingat
var
;
vars
CautionsSkrift
ock
nu
presenterades
.
§
6
.

Sedan
innehavarna
av
Skräptorphemmanet
,
levererat
till
Fattighuset
sin
spannmjöls
Ränta
för
förra
året
,
men
icke
penningskatten
;
bestigande
sig
till
9
dal
.
31
Va
öre
kmt
,
förfrågade
sig
Kyrkoherden
:
om
han
skulle
lagligen
utsöka
dessa
penningar
?

Tillsades
Församlingen
,
av
Nämndemannen
,
å
Landsman
Hinsings
vägnar
,
att
forderligast
reparera
sina
Brolotter
,
vid
den
av
vattufloden
fördärvande
Forssiöbronn
.
§
32
.

Lät
Kyrkoherden
Församlingen
veta
det
han
,
strax
efter
den
nyligen
timade
Hemming
Swänssons
död
låtit
uti
Fattighuset
igenom
sin
Adjunkt
Herr
)
öjerstedt
och
bägge
Fattigfogdarna
,
vederbörligen
inventera
all
dess
kvarlåtenskap
,
samt
att
efter
bemälte
Hamming
då
funnits
213
dr
28
.
/
.

Begärde
Pastor
,
att
Församlingen
ville
sig
utlåta
om
avlidne
Nummer
soldaten
Malmquists
dotter
,
som
nu
igenom
kyrkoherdens
Kristliga
försorg
lärt
läsa
så
mycket
,
som
hon
i
sin
sinnens
svaghet
fatta
kan
,
längre
skulle
vara
i
fattighuset
Församlingen
till
last
och
tunga
,
samt
om
någon
av
närvarande
Socknens
invånare
kunde
och
visste
giva
förslag
på
någon
tjänlig
tjänst
för
henne
;
Per
Andersson
uti
Remmerö
med
flera
,
intygade
,
det
de
ej
det
göra
kunde
,
särdeles
som
Flickan
efter
deras
mening
ännu
ej
skulle
kunna
någon
tjänst
förestå
,
samt
att
väl
vore
om
någon
av
anhöriga
här
efter
ville
henne
vårda
;
Varpå
slikt
blev
belovat
,
att
Flickan
skulle
igenom
någon
viss
beskedlig
Karl
,
förmedelst
Pastoris
försorg
,
föras
till
sin
Faster
uti
Wingåkers
östra
Församling
som
barnlös
är
,
och
stå
under
dess
vård
intill
dess
hon
denna
sin
Brorsdotter
ställa
kan
i
tjänst
som
Flickan
kan
vara
belåten
vid
.
§
10
.

Herr
Löjtnanten
Lidstrand
,
såsom
mesta
rösterna
ägande
i
Församlingen
,
berättade
sig
denna
saken
ännu
ej
ha
nog
övervägt
:

Sedan
Församlingen
berättat
hade
,
att
den
på
sista
Valborgmässosockenstämman
,
av
Påhlstorpa
rota
föreslagna
skomakaren
ifrån
Juhlita
,
på
den
orten
fått
lägenhet
,
och
därför
icke
hit
anlänt
,
frågade
Pastor
om
Lars
Gustafsson
måg
uti
Porten
,
efter
det
slut
,
som
träffat
blev
på
sist
hållna
Valborgsmässo
Sockenstämman
,
så
hade
betjänt
Församlingens
invånare
uti
Kåhlmån
,
att
de
med
hans
Skoarbete
kunde
vara
förnöjda
.

Vederbörande
svarade
;
att
icke
någon
med
skäl
uppå
hans
arbete
kunde
ha
till
att
klandra
utan
ville
gärna
ha
denna
mannen
här
efter
för
sin
hantverkare
.

Ville
Pastor
ha
föravskedade
Nummer
Soldaten
Lars
Norman
varnat
,
att
ej
bruka
någon
lärogosse
vid
sitt
skräddarehantverk
,
Församlingens
gärningsmän
,
emot
förordningen
,
till
förfång
.

Efter
saligt
avlidne
Kyrkovärden
Per
Persson
i
Stensiö
,
som
i
20
år
sysslan
haft
vid
Kyrkan
,
och
densamma
med
all
trohet
förvaltat
,
blev
Nämndemannen
Nils
Nilsson
uti
Remna
,
med
Församlingens
enhälliga
samtycke
,
till
Kyrkovärd
antagen
.
§
10
.

Herr
Löjtnanten
Lidstrand
tyckte
bäst
vara
detta
stycket
att
omlaga
med
grovt
ör
som
kunde
tagas
ifrån
hemmanet
Väggen
uppå
Monn
;
vartill
även
den
övriga
Församlingen
samtyckte
,
slutandes
att
de
närmst
intill
Kyrkan
boende
skola
köra
tvenne
parlass
för
ett
dagsverke
.
§
17
.

För
denna
skull
begärde
Pastor
Församlingens
utlåtelse
över
detta
Lars
Perssons
egenvilliga
förhållande
.

Gav
Pastor
vid
handen
,
att
han
efter
överenskommande
på
sistlidna
Sockenstämma
;
ej
kunnat
låta
göra
nytt
golv
uti
Sockenstugan
,
och
det
av
brist
på
tjänligt
tegel
;
men
försäkrade
framdeles
att
vilja
draga
behörig
försorg
,
huru
bemälte
golv
med
tjänliga
tegelstenar
måtte
lagt
varda
.
§
8
.

När
detta
så
var
belovat
förklarade
sig
Sockenskräddarna
Sven
Svensson
ej
kunna
vara
nöjd
med
denna
taxa
;
blev
därför
föravskedad
,
och
kvitt
de
förmåner
,
som
han
genom
sitt
hantverk
i
denna
församlingen
ägt
och
haft
'
.
§
10
.

Desslikes
berättade
Komministern
Georg
Netzelius
det
han
av
sin
dräng
fått
höra
,
att
denna
gosse
sistlidna
andra
Bönedag
försummat
gudstjänsten
,
fast
än
han
varit
vid
kyrkan
,
som
Brodern
till
Komministerns
dräng
,
föravskedade
Nummersoldaten
Lars
Norman
för
drängen
berättat
.

Fjärde
Bönedagen
ingen
såsom
absens
annoterad
;
med
allvarsam
tillsägelse
,
att
dessa
skola
äntligen
igenom
verifikationer
bevisa
,
antingen
att
de
varit
vid
Gudstjänsterna
på
dessa
Bönedagar
uti
andra
kyrkor
i
grannskapet
eller
ock
att
de
haft
giltiga
orsaker
till
deras
hemma
blivande
,
och
det
åtta
dagar
för
instundande
hösteting
,
så
skönt
de
ville
undvika
att
bli
lagförda
.
§
21
.

Så
lovade
även
Pastor
att
skänka
henne
litet
ull
till
kläder
åt
det
fattiga
barnet
.
§
27
.

Emot
alla
dessa
tydliga
räkningar
hade
ingen
något
att
påminna
utan
erkändes
alltsammans
ha
sin
riktighet
.
§
3
.

Beviljade
Församlingen
Lars
Pärssons
hustru
uti
Rössnebo
(
=
Rosselbo
)
,
Fattigdel
,
ibland
)
allmosehjonen
,
utom
Hospitalet
,
i
anseende
till
dess
blindhet
och
stora
Sjukdom
.

Men
detta
målet
blev
till
ett
annat
tillfälle
uppskjutet
.
§
10
.

Förmanades
ock
Ämbetsmännen
,
vilka
nu
även
tillstädes
var
,
att
ställa
sig
denna
Församlingens
överenskommelse
,
till
behörig
efterrättelse
,
och
för
all
ting
göra
sitt
arbete
,
alldenstund
den
så
tillräcklig
arbetslön
beviljad
är
,
med
den
tro
och
uppriktighet
,
som
de
bäst
försvara
kunde
.

§
.
uti
sisthållna
Mickelsmässo-Sockenstugo-Protokoll
berättade
Herr
Probsten
,
det
Kamreren
vid
Claestorp
Herr
Pehr
Sundling
,
efter
församlingens
gottfinnande
varit
här
ock
,
förrän
Orgel-nisten
Pehr
Oxelberg
flyttat
hädan
till
Arboga
Stad
,
inventerat
ifrån
honom
orgelverket
härstädes
,
som
befanns
riktigt
,
varöver
även
bemälte
Herr
Kamreren
givit
sitt
skriftliga
vittnesbörd
.
§
13
.

Vid
samma
tillfälle
befalldes
Walla
Rotes
Sexman
,
nämligen
Lars
Larson
i
St.
Fräntorp
,
att
gå
till
Tohlgiölet
,
innan
Brita
flyttar
in
i
fattighuset
,
och
noga
se
efter
vilka
saker
hon
har
med
sig
,
som
böra
efter
lag
och
Tiggareordningen
komma
fattighuset
till
tjänst
efter
hennes
död
.

Framkallades
unga
Tjänstedrängen
Gustaf
Ersson
uti
Harstorp
,
tillika
med
drängen
Pehr
Pehrsson
i
Walla
,
av
vilka
den
förre
allvarsamt
förehölls
det
grova
ofog
han
emot
den
senare
förövat
,
samt
huru
mera
bestialiskt
,
än
naturligt
,
han
någon
tid
tillförende
,
under
deras
Hoparbete
honom
hanterat
,
med
flera
föreställningar
,
för
att
honom
erinra
dess
vanart
;
Påmindes
jämväl
,
att
ändock
Respektive
Herrskapet
på
Ericsberg
,
av
högtberömlig
nit
för
ordning
och
Kristlig
sedighet
ibland
sitt
folk
,
honom
behörigen
korrigerat
m.m.
borde
han
icke
desto
mindre
nu
,
både
bedja
Församlingen
om
förlåtelse
,
som
han
,
jämte
den
rättfärdige
Guden
,
igenom
sin
odygd
förtörnat
och
förargat
,
såsom
ock
till
Pehr
Pehrsson
betala
den
förlikning
,
högbemälda
Herrskap
honom
med
all
rätt
pålagt
,
innan
han
må
tänka
sig
admitteras
till
den
Heliga
Nattvarden
,
m.m.
Det
förra
gjorde
Gustaf
strax
,
bekännande
sig
ha
rätt
illa
gjort
,
och
det
senare
lovade
Gustafs
fader
,
innan
aftonen
erlägga
och
betala
.

Avsade
sig
Sexmans
Sysslan
Pehr
Pehrsson
i
Högen
,
Lars
Larsson
i
St.
Fräntorp
och
Eric
Persson
i
Remmarö
,
och
uti
deras
ställen
förordnades
Pehr
Hansson
uti
Brenäs
,
Anders
Olson
i
Åbohl
och
Olof
Pehrsson
i
Klicksta
.
§
24
.

Till
Lars
Olsons
fattiga
moder
uti
Kålstugan
,
lovade
ock
Församlingen
någon
hjälp
,
i
varande
svåra
tid
,
så
mycket
Fattigkassan
kunde
tillåta
.
§
25
.

Anmodades
Föreståndarna
för
Socken
Magasinet
,
att
vid
nästa
Intäkten
,
av
den
i
Somras
utlånade
Spannmålen
,
vara
,
efter
vanligheten
,
behjälpliga
,
som
utlovades
.
$
11
.

Som
ett
parti
Sågbockar
och
Plankstycken
är
vid
Kyrkan
övriga
,
efter
det
till
SockenMagasinet
Sågade
Timmer
,
vilka
på
intet
sätt
kunna
för
Kyrkans
behov
employeras
Så
biföll
Församlingen
det
förslaget
,
att
på
någon
lätthelgedag
i
höst
,
besagda
Persedlar
kunde
för
kyrkans
räkning
förauktioneras
.
§
14
.

Andra
i
Församlingen
invände
,
att
deras
gärningsmän
har
tyskt
Skoarbete
ofta
förhänder
,
varigenom
sker
,
att
vederbörande
Rotars
Åbor
icke
kunna
betjänas
som
de
borde
;
Herr
Probsten
utlät
sig
häröver
,
att
detta
målet
icke
till
denna
,
utan
nästkommande
Mickels
MässoSockenStämman
hörde
;
I
vilket
avseende
,
det
ock
blev
denna
resan
uppskjutet
,
med
erinring
,
att
förenämnda
osed
borde
avskaffas
,
och
vederbörande
gärningsmän
allenast
hålla
sig
vid
det
svenska
Skoarbetet
till
Rotarnas
så
mycket
bättre
betjänande
.
§
7
.

Församlingen
tog
fuller
detta
ärendet
uti
vederbörligt
övervägande
;
man
fann
sig
icke
befogad
att
utsätta
någon
viss
vedergällning
Johan
Bengtson
till
förmån
för
sitt
omak
med
dessa
foror
årligen
,
utan
tyckte
rådligast
vara
,
att
uppskjuta
målet
till
ett
annat
tjänligt
tillfälle
.
§
17
.

November
samma
år
,
utsynt
till
SockenMagasinet
,
till
antalet
400
stycken
,
var
allenast
till
Kyrkan
framskaffade
,
161
Såg
och
Timmerstockar
tillsammans
räknade
,
så
att
ännu
återstå
,
174
Såg
och
65
Timmerstockar
,
tillsammans
239
stycken
,
vilka
den
19
November
1761
blev
av
den
nuvarande
Skogvaktaren
Johan
Öberg
,
utsynade
.

Att
man
icke
annat
hört
och
vet
,
än
allt
som
är
under
främsta
valvet
,
varest
ock
ifrån
de
äldsta
tider
tillbaka
,
de
ifrån
Djula
avlidna
,
finnas
begravna
.
§
21
.

Begärandes
därjämte
,
att
Pastor
ville
,
vid
tillfälle
,
med
Högvälborne
Herrn
Hovmarskalken
,
om
de
förmälda
revor
på
Hörnen
av
Gaveln
,
och
deras
botande
överlägga
,
och
låta
sedermera
,
Herr
Löjtnanten
därav
del
få
.
§
26
.

Och
påmindes
:
att
sådant
,
jämte
dagsverken
,
borde
ske
med
Församlingens
Kostnad
och
icke
Kyrkans
,
vartill
samtycktes
i
proportion
på
hemmanen
.
§
14
.

Välborna
Fru
Lagmanskan
Rosenstam
på
Wärhulta
,
begärde
några
flera
,
av
Församlingen
,
underskrift
,
jämte
Kyrkoherdens
,
på
Cautionen
för
Frälsehemmanet
Banninge
,
som
av
Orgelnisten
arrenderas
;
vilket
ock
nu
skedde
.
§
18
.

Gav
Sockenskomakaren
Lars
Larsson
i
Harbacken
tillkänna
,
att
han
icke
längre
än
till
nästa
Michaelii
,
kan
tjäna
församlingen
med
sitt
arbete
.
§
20
.

Martii
sistledne
,
som
även
nu
upplästes
,
innan
nästa
mantalsskrivning
,
göra
sig
noga
underrättade
om
både
gamla
och
unga
i
alla
hushållen
,
på
det
Hans
Kungl.
Majts
Nådiga
befallning
,
i
all
måtto
må
efterlevas
;
och
lovade
Pastor
att
av
Predikstolen
,
när
rätta
tiden
i
höst
,
vill
Gud
,
infaller
,
därom
påminna
.
§
22
.

Som
mantalsskrivningen
snart
tillstundar
,
frågades
:
om
något
ombyte
sker
med
Socknens
gärningsmän
?

Vad
en
gång
,
med
Församlingens
allmänna
gottfinnande
skett
,
borde
nu
icke
dragas
till
Exempel
,
emedan
det
både
är
emot
alla
Församlingars
praxis
,
såsom
ock
vet
man
ingen
förordning
diktera
,
att
de
reparationer
som
ske
utom
Bogårdsmuren
,
bör
ske
för
Kyrkans
kostnad
.

Men
som
det
nu
varande
Fattighus
förrådet
sådant
icke
,
utan
brist
och
saknad
för
de
andra
,
kunde
,
lovades
henne
någon
hjälp
ifrån
Prästgården
.
§
14
.

Anmodades
,
av
Församlingen
,
Sockenskräddaren
Petter
Olofsson
,
att
i
höst
uti
lära
antaga
den
fader
och
moderlösa
gossen
Eric
Olson
,
vars
moder
,
Ingeborg
Hansdotter
,
nyligen
förut
i
Fattighuset
avlidit
,
vilket
han
ock
lovade
,
så
vida
han
ville
sig
beskedligen
skicka
och
förhålla
.
§
3
.

I
avseende
därtill
blev
Lars
Carlsson
i
Foglö
och
Johan
Bengtsson
i
Wrå
,
föreslagna
;
då
igenom
lättande
,
Lars
Carlsson
,
förordnades
till
Kyrkovärd
.
§
9
.

Som
även
man
förmärkt
,
att
drängar
och
Pigor
nu
mera
förgätit
det
förbud
och
vite
,
som
Församlingen
sig
emellan
fastställt
,
så
väl
på
Mickelsmässo
Socken
Stämman
den
)
29
.

Så
upplästes
icke
allenast
förenämnda
Socken
Stämmo
Protokoll
,
utan
förekallades
ock
tjänstedrängen
Jonas
Eliason
uti
Kårtorp
,
och
tilltalades
allvarsamt
,
tillika
med
Nummer
Soldaten
Malmstedt
,
den
förre
för
det
han
nyligen
tillförende
,
under
nattvardsgången
understått
sig
med
blå
knappar
i
kyrkan
komma
;
den
senare
för
det
han
,
efter
berättelse
,
har
en
sådan
Rock
förfärdigat
.

Uppräknades
de
som
restera
med
den
vanliga
Veden
,
för
nästlidna
vintertid
till
Fattighuset
,
och
tillsades
Sexmännen
,
att
tillsäga
vederbörande
det
de
vid
förr
utsatta
vitet
,
med
första
sin
skyldighet
fullgöra
.
§
18
.

Församlingen
icke
vidare
kunde
sig
med
målet
befatta
.
§
6
.

Som
ock
det
blivit
av
Murmästaren
österberg
,
tillkännagivet
,
under
det
han
med
kyrkodagsverkarna
på
nya
Koret
var
sysslosatt
,
det
mera
nämnda
drängar
Anders
Andersson
)
och
Pehr
Olofsson
,
efter
utståndet
straff
den
)
4
i
denna
månad
,
har
på
en
vagn
åkandes
förbi
kyrkan
,
skrikit
och
ropat
,
samt
eljest
oanständigt
sig
betett
:

Berättade
även
Pehr
Nilsson
uti
Harstorp
,
på
tillfrågan
om
samma
ärende
,
att
hans
Son
Anders
hade
sig
målet
bäst
bekant
.
§
9
.

Vad
han
på
dessa
4
vittnens
enhälliga
utlåtande
,
och
dem
han
icke
gittat
jäva
,
hade
att
svara
?

Lars
Larssons
hustru
i
Opsala
,
som
varit
anmodad
att
besiktiga
barnet
,
berättade
:
att
barnet
varit
litet
blått
på
högra
kindbenet
,
och
haft
en
liten
rödstrimma
neder
åt
näsan
;
Eljest
hade
hon
ingen
åkomma
skönja
kunnat
.
§
3
.

Om
hon
vårdat
och
älskat
sitt
barn
,
eller
om
det
vanskötts
av
henne
,
m.m.
?
Vartill
svarades
:
att
ingen
visste
annat
än
det
som
beskedligt
var
.
§
4
.

§
.
13
.
samt
den
i
alla
Församlingar
lovligen
)
vedertagna
plägesed
,
nästkommande
Söndag
sätta
sig
uti
den
nedersta
Kyrkobänken
,
och
med
Församlingen
troligen
förena
sina
böner
till
den
Barmhärtiga
Guden
,
efter
det
Formulär
,
som
uti
Hand
Boken
beskrivet
finns
,
och
sedermera
om
Gud
Henne
med
någon
livsfrukt
vidare
välsigna
täcktes
,
lära
sig
vakta
för
vårdslöshet
m.m.
Så
vara
hänt
,
intygar
på
Församlingens
vägnar
,
J
.
Dalenius
P
.
&
Pr.p.t.l
.

Ehuru
Boström
emot
detta
vittnet
;
intet
hade
att
invända
,
framfor
han
icke
desto
mindre
uti
sina
förra
obetänkta
utlåtelser
,
oaktade
alla
till
honom
skedde
allvarsamma
varningar
,
sägandes
:

Juni
,
hölls
,
efter
2
dagars
förut
skedd
kungörelse
av
Predikstolen
,
Alman
Valborgsmässo
Sockenstämma
,
i
närvaro
av
Församlingens
respektive
Herrskapers
Betjänter
,
Socknens
äldsta
och
Sexmän
,
med
)
flera
)
då
följande
avhandlades
.

Rekommenderade
församlingen
,
efter
följande
Hus
fattiga
,
någon
hjälp
av
FattigKassan
,
såsom
Pehr
Pehrsson
i
Sandbäckstufwan
,
9:dr
.

Tackade
man
församlingens
invånare
,
för
dess
enhällighet
,
att
uti
förvekne
Höst
och
Vinter
,
riktigt
betala
det
vanliga
matskottet
av
veden
till
fattighuset
,
och
uppräknades
de
med
ved
resterande
,
Stora
)
och
Lilla
)
Fräntorp
,
Gafwelen
,
Sjöstufwan
,
Tohlgölet
,
Tohltorp
,
Elgsjötorp
,
Källstufwan
,
Olofstorp
,
Sundstufwan
och
Anders
Andersson
i
Remmerö
,
allt
för
1766
,
men
med
det
vanliga
matskottet
,
resterande
allenast
Sundstorp
.

Utfästande
sig
Sexmännen
,
att
vid
nästa
Vinterföre
,
sådant
infordra
.
§
11
.

Om
det
icke
vore
dess
vilje
,
att
för
Fattigmedlen
någon
Fattigbössa
vid
Stensjö
upprättades
,
varav
man
kunde
något
vid
vissa
tillfällen
,
så
under
påstående
Ting
,
som
av
resande
,
förvänta
,
alldenstund
igenom
Utdrag
av
Protokollet
,
den
)
3
November
1767
,
/
:
som
nu
även
upplästes
,
/
Härads
Rätten
därtill
sitt
bifall
lämnat
?

Huruvida
Församlingen
ville
till
efterlevnad
antaga
den
av
Högvälborne
Herr
Greven
,
Kommendören
och
Landshövdingen
Nils
Bjelke
,
utgivna
ByOrdningen
tillika
med
den
av
honom
författade
Underrättelsen
,
huru
man
i
missväxts
år
,
med
ringa
möda
och
särdeles
Hö
och
SädesBesparing
,
kan
framföda
,
drag
och
andra
Kreatur
.

I
anledning
därav
utbad
man
sig
Församlingens
benägna
utlåtande
,
på
vad
sätt
både
denna
fordran
måtte
betalas
,
såsom
ock
om
det
kunde
tillåtas
,
att
någon
privat
person
i
församlingen
,
finge
för
sin
räkning
insätta
några
Tunnor
,
emot
IV2
Kappars
betalning
av
Räntan
,
till
Magasinet
årligen
?

Första
resan
sistledne
midsommarafton
,
och
sedermera
flera
resor
,
men
sista
gången
nästförut
gående
Torsdag
,
eller
den
)
20
Juli
,
då
hon
ock
skall
ha
kört
upp
hennes
kor
ifrån
mossen
.
§
3
.

Upplästes
Boken
och
Fattig
Kassans
utestående
fordringar
och
underskrevs
.

Till
slut
bad
han
om
förlåtelse
och
lovade
förbättring
.
§
20
.

Gubben
i
Ändebol
kunde
icke
intagas
i
fattigstugan
,
helst
intet
rum
nu
var
ledigt
.
§
29
.

Vartill
Herr
Inspektorn
täcktes
sitt
bifall
och
löfte
lämna
.

Församlingens
förnäma
Patron
lät
giva
tillkänna
,
att
han
förordnat
unga
Herr
lan
Eric
Oxelberg
till
Orgelnistsysslans
bestridande
härstädes
tills
vidare
,
och
att
bemälte
Oxelberg
äga
uppbära
därför
så
stor
Spannmålslön
av
församl:n
,
som
hans
företrädare
njutit
.
6:o
.

Pastor
har
anmärkt
,
hur
några
äkta
makar
följa
varandra
fram
till
den
Hel
.
nattvardens
undfående
,
men
de
flesta
icke
så
,
varigenom
händer
,
att
gifta
och
ogifta
,
gamla
och
unga
,
blanda
sig
om
vartannat
,
vilket
icke
utmärker
den
ordning
och
skick
vid
nattvardsgången
,
som
nästan
överallt
i
alla
församlingar
i
Riket
är
brukligt
.

Församlingen
tog
detta
mål
i
övervägande
och
beslöt
enhälligt
,
att
alla
nattvardsgäster
skola
hädanefter
och
allt
framgent
följa
och
iakttaga
denna
ordning
,
som
aldrig
skall
ändras
och
består
däruti
,
att
vid
den
h
.
nattvardens
anammande
skola
först
alla
gifta
män
,
var
och
en
med
sin
hustru
,
falla
på
knä
bredvid
varandra
,
sedan
framträda
alla
ogifta
söner
och
drängar
och
sist
framkomma
alla
ogifta
döttrar
och
pigor
.

Vad
änklingar
och
änkor
angår
,
så
kunna
de
följa
med
de
gifta
.

Församlingen
tyckte
,
att
detta
priset
var
ganska
billigt
,
och
beslöt
,
att
räkningen
skulle
nu
betalas
.
§
20
.

På
begäran
beviljades
Sexmannen
i
Rcmna
avsked
,
och
antog
församlingen
nu
till
Sexman
i
kyrkoroten
Sockenmannen
Lars
Larsson
i
Stensjö
.
§
25
.

Församl:n
trodde
,
att
om
Pastor
på
predikstolen
föreställde
detta
genom
ett
lämpligt
tal
,
så
skulle
de
i
denna
saken
brottsliga
taga
sig
till
vara
och
visa
lydnad
.

Och
beträffande
den
gamla
byggningen
,
önskade
jag
att
den
obrukbara
delen
därav
kunde
under
byggnaden
rivas
,
så
att
åtminstone
bräderna
uti
tak
och
bölning
fingo
användas
vid
den
nya
byggnaden
,
såsom
förmånligast
för
församl:n
,
ty
det
förstås
av
sig
själv
,
att
den
delen
,
som
nu
av
Pastor
bebos
,
ej
kan
föryttras
el:r
till
församlingens
hjälp
användas
,
innan
nya
huset
blir
bebott
.

Sammaledes
förhålla
det
sig
med
dörrarna
,
när
Psalmen
efter
predikan
börjas
,
så
att
ingen
får
gå
ur
kyrkan
,
förrän
allt
är
slutat
.

Häröver
beslöts
,
att
om
han
icke
tjänar
här
i
Socknen
,
utan
sitter
blott
i
hus
,
borde
han
tillsägas
,
att
begiva
sig
till
sin
ort
igen
,
men
i
annan
händelse
icke
.
§
19
.

Jag
är
genast
färdig
att
för
mina
underhavande
i
socknen
uti
denna
del
följa
lagens
bokstav
,
varigenom
jag
fredas
ifrån
vidare
ändring
av
vad
en
gång
blivit
beslutat
.

Sedan
alla
resp
.
jordägare
genom
sina
fullmäktige
och
alla
jordbönderna
själva
församlat
sig
i
Sockenstugan
,
att
överlägga
om
antagandet
av
den
på
10
år
av
Kungl
.

Alla
närvarande
förmenade
sig
ha
inhämtat
tillräcklig
.
kunskap
härom
.

Fjärdingsmannen
frågade
dem
härvid
,
vad
de
hade
mot
hans
Kungl.
Maj:ts
nådiga
anbud
?

Carl
Andersson
i
Kerstinboda
förehölls
och
tillsades
allvarsamt
att
avstå
med
sitt
buller
i
Kyrkan
och
med
sin
obeskedlighet
i
de
hus
,
han
besöker
.

Som
man
tyckte
,
att
penningsammanskottet
allenast
av
3
rotar
till
ljus
om
Julottan
blev
för
litet
;
så
vart
beslutat
,
att
det
årligen
skulle
utgöras
av
4
rotar
.

Upplästes
,
godkändes
och
underskrevs
,
såväl
de
sist
hållna
protokollen
,
som
ock
räkenskaperna
över
Kyrko
och
fattigkassorna
.
§
2
.

Och
som
denna
Psalm
sjunges
vid
början
av
varje
kommunion
,
då
orgelverket
icke
nyttjas
,
så
förmenade
Pastor
,
att
församl:n
kan
då
bäst
höra
och
akta
på
,
hur
organisten
sjunger
och
vid
vilka
ord
han
håller
litet
upp
,
och
således
därav
lära
sig
sjunga
rätt
.
§
7
.

S
.
pag.
520
,
§
2.22
)
4:o
Beviljades
gamle
Jon
i
Löfåsen
full
fattigdel
eller
i
l:sta
klassen
,
men
kommer
att
ha
husrum
hos
sin
Son
.

Han
svarade
,
att
på
auktion
vid
Julfors
hade
ett
ganska
oskickat
väsende
förelupit
,
men
för
sina
göromål
skull
hade
han
icke
haft
tillfälle
att
själv
kunna
se
,
vilka
de
varit
,
som
det
utövat
.

Lind
tillkännagav
församl:s
Herr
Patroni
vilja
,
att
nästa
vår
skola
alla
stolar
i
kyrkan
nedtagas
,
golvet
över
allt
planeras
och
nya
stolar
åter
insättas
.

C
.
h
.
Uggla
.
"
Som
ändamålet
med
besvarandet
av
föreskrivna
frågor
,
skulle
vara
,
att
bereda
Herr
Kammarherrens
yttrande
i
den
redan
i
Sockenstämma
av
St.
Malms
församl
.
avgjorda
frågan
om
tomma
Magasinshusets
försäljande
,
kunde
sådant
skäligen
synas
överflödigt
;
men
då
Herr
Kammarherrens
önskan
därjämte
tymedelst
kan
tillfredsställas
,
anser
jag
för
ett
nöje
,
att
därom
punktvis
lämna
följande
svar
:
l:o
.

Hur
vissa
inrättningar
och
behov
ej
där
kunna
äga
rum
,
känner
H:r
Kammarherren
förut
,
som
behagade
föra
sig
till
minnes
,
att
till
exempel
kroginrättningar
på
kyrkovallen
ej
är
tillåtna
.

Linds
uti
sista
Sockenstämma
anmälda
utlåtande
,
att
med
Magasins
husets
försäljande
upskjutas
tills
efter
andetiden
,
är
jag
så
mycket
mer
tillfreds
,
som
jag
nu
avreser
från
orten
,
men
,
vill
Gud
,
i
början
av
Sept
.
tänker
vara
återkommen
,
då
om
auktionsdagen
får
samrådas
.

På
stenen
var
samma
personer
,
fast
i
större
skapnad
,
uthuggna
,
som
stå
avmålade
på
den
tavlan
,
vilken
hänger
på
muren
där
bredvid
,
samt
med
bokstäver
omkring
.

Djula
ägares
rätt
till
gamla
koret
i
St.
Malms
kyrka
har
förut
aldrig
blivit
bestridd
,
varför
jag
så
mycket
mindre
väntat
mig
ett
så
ovänligt
steg
av
Ericsbergs
ägare
.

Och
bör
detta
Häradsrättens
förbud
till
vederbörl
.
efterrättelse
offentl
.
kungöras
,
på
det
ingen
okunnighet
därav
,
om
det
på
något
sätt
överträdas
skulle
,
förebäras
och
invändas
må
.

Åliggandes
jämväl
H:r
Hovauditören
Ehrenfelt
,
att
vid
nästa
ting
inkomma
,
om
han
något
vid
stolläggningen
har
att
andraga
eller
vara
sin
talan
förlustig
.

Uti
Herr
Kammarherren
Uggla
äger
församl:n
en
kunnig
ledamot
,
som
säkert
gör
sig
ett
nöje
att
gagna
och
vars
tid
även
torde
lämna
honom
ett
därtill
gott
och
tjänligt
rådrum
.

Herr
Patronus
tillsade
,
att
kyrkan
med
det
första
skall
göra
avbetalning
på
denna
skuld
,
allenast
så
mycket
behållas
kvar
i
kassan
,
som
fordras
till
Kommunion
vins
inköpande
och
andra
nödiga
utgifters
bestridande
,
skänkande
Herr
Patronus
efter
Intressen
på
skulden
.

Prosten
nämnde
,
att
ett
rum
vore
ledigt
i
fattigstugan
och
även
en
full
fattigdel
utom
,
samt
för
en
person
i
2dra
klassen
.

Herr
Patronus
täcktes
svara
,
att
om
bodarna
var
bristfälliga
för
7
år
sedan
,
vad
skola
de
då
nu
icke
vara
,
begärde
få
höra
ur
husesyns
Dokumentet
,
som
nu
var
tillhands
,
vad
Synerätten
prövat
åtgå
till
dessa
Bodars
byggande
,
och
biföll
nybyggnaden
,
med
det
påstående
,
att
den
bör
auktioneras
till
den
minst
bjudande
.

Maneck
,
Pr
.
et
P
.
Uppläst
och
till
alla
delar
erkännes
av
Gerhard
Lind
Pehr
Pehrsson
i
Brenäs
Efter
fullmakt
nämndeman
Olof
Pärsson
i
Banninge
Erik
Andersson
i
Walla
Kyrkovärdar
Olof
Erickson
i
Gersnäs
Lars
Jönsson
i
Stensiö
Lars
Jonsson
Sexmän
Erick
Persson
i
Remrö
Eric
Ersson
i
Remrödstorp
Benet
Pehrsson
i
Remrö
År
1790
den
17
Oktober
.
inträdde
församl:s
Invånare
uti
Sockenstugan
,
att
justera
det
vid
sista
allmänna
Mickelsmässo
Sockenstämman
hållna
protokoll
.
§
1
.

Min
Fullmäktig
är
alltså
berättigad
,
att
vid
den
sammankomst
,
som
i
dag
hålles
,
så
uppföra
sig
,
som
om
jag
själv
vore
närvarande
,
samt
i
skrift
el:r
tal
anföra
,
rätta
,
påminna
el:r
tillägga
,
vad
han
finner
till
saken
hörande
och
till
mina
rättigheters
försvar
ländande
,
vilket
jag
för
gott
anser
.

H:r
Mag:r
Duvser
sade
,
att
ingen
måtte
kunna
åtaga
sig
det
för
sålitet
.

H:r
Patronus
svarade
:
ja
,
jag
erkänner
det
till
alla
delar
.
§
6
.

Kvittensen
var
av
detta
innehåll
:

Till
yttermera
visso
varder
detta
kvittens
av
mig
egenhändigt
underskrivet
och
med
mitt
vanliga
signet
bekräftat
,
som
skedde
i
Stockholm
d
.
12
Maj
1795
.

Jacobson
sigill
I
anledning
härav
framgav
Herr
Bruksinsp
.
Lind
till
uppläsande
en
lista
,
underskriven
av
Ericsbergs
Possessor
Välb.
Herr
David
Gotthard
Hildebrand
,
på
15
fattiga
personer
,
som
välbemälda
Herre
behagat
nämna
till
åtnjutande
av
de
lOOde
Rdr
,
vilka
emellan
dem
så
utdelas
skulle
,
att
vardera
fick
6
Rdr
32
s
.
-
Dessa
lOOde
Rdr
blev
ock
nu
genom
Bruksinsp
.
Lind
till
Prosten
och
de
2ne
fattigkassans
föreståndare
överlämnade
,
som
dessa
pgr
till
de
utnämnde
15
fattiga
utdela
skulle
och
på
vilken
summa
de
nu
kvittens
gav
.
-
Fattigkassans
föreståndare
fann
för
gott
,
att
till
dessa
fattiga
nu
utdela
endast
halva
summan
och
den
andra
hälften
fram
åt
Olofsmässan
,
för
att
förmå
dem
,
att
desto
bättre
med
denna
stora
nådesgåvan
hushålla
och
vartill
de
även
nu
föreställningar
undfick
.
§
3
.

Varför
nu
beslöts
,
att
vart
matlag
hädanefter
ger
därtill
1
s.
,
och
skulle
något
överbliva
av
dessa
pgr
,
sedan
18
r
talg
är
uppköpta
,
så
tillfaller
det
kyrkokassan
.
§
10
.

Sedan
församlingen
sport
,
att
v
.
Häradsdomaren
Pehr
Pehrsson
i
Brenäs
vid
instundande
höstting
i
Stensjö
tänker
begära
avsked
,
och
som
en
nämndeman
alltid
varit
i
denna
socken
boende
,
den
därstädse
varit
sysselsatt
med
de
mål
,
hans
kallelse
honom
ålagt
;
så
fann
församlingens
invånare
nödigt
,
att
i
denna
blivande
ledigheten
i
dag
utse
och
föreslå
3ne
ärliga
och
förståndiga
män
av
sina
medlemmar
,
samt
stannade
i
det
beslut
,
att
på
nämndemans
förslag
uppföra
frälse
bönderna
Pehr
Ersson
i
Stensjö
,
Lars
Nilsson
i
Stensjö
och
Olof
Ersson
i
Fogelö
,
åstundades
,
att
detta
förslag
medelst
utdrag
av
protokollet
hos
välborne
Herr
Häradshövdingen
å
hösttinget
med
Oppunda
härad
måtte
anmälas
,
under
avvaktan
av
dess
gunstiga
utnämnande
.

Upplästes
,
erkändes
och
underskrevs
så
väl
sisthållna
protokoll
,
som
ock
räkenskaperna
över
Kyrko
och
fattigkassorna
.
§
2
.

Jan
Jonsson
i
Mokällan
blev
på
sin
begäran
från
sockenskomakarverket
entledigad
.
§
8
.

Martii
,
i
anledning
av
Häradshövding
välborne
Herr
v
.
Jacobsons
kungörelse
,
att
Oppunda
Härads
boer
komma
att
inställa
sig
d
.
12
nästa
Martii
i
Stensjö
,
till
att
syna
det
bristfälliga
Tingshuset
och
överenskomma
om
dess
förbättrande
,
inkallades
denna
församlingens
invånare
,
att
utnämna
sin
fullmäktig
vid
ovannämnde
mål
,
och
föll
de
med
sitt
förtroende
på
v
.
Notarien
i
Kungl.
Svea
hovrätt
,
ädel
och
högaktad
Herr
Anders
Lindblad
,
att
vara
deras
befullmäktigade
ombud
,
förklarande
sig
nöjda
med
vad
Herr
Notarien
härutinnan
lagl
.
(
igen
)
gör
och
låter
.

April
blev
Extra
Sockenstämma
hållen
med
St.
Malms
församling
)
efter
föregången
pålysning
.

Summan
skulle
utdelas
i
2ne
terminer
,
såsom
tillförene
skett
.
4o
.

Detta
ärendet
åtog
sig
nu
org
.
Humla
och
varvid
församl
.
ålade
honom
1
Rdrs
böter
för
var
gång
han
försummar
verkställa
någon
gravöppning
,
av
vilka
böter
gravöppningen
då
av
en
annan
göres
och
överskottet
tillfaller
fattigkassan
.

Sexman
i
Prästorp
anförde
,
att
en
nyl
.
gift
hustru
från
Lerbo
,
som
förr
tjänat
i
Valla
och
vars
man
nu
tagit
tjänst
i
Sköldinge
,
hade
flyttat
till
Sandstug
.

Av
hkn
(
vilken
)
anledning
de
,
efter
kungörelse
från
predikstolen
,
nu
tillstädes
kom
,
och
,
underrättade
om
ändamålet
med
deras
sammankallande
,
instämde
enhälleligen
däri
,
att
vända
sig
till
Länets
Styresman
,
för
att
i
ödmjukhet
utbedja
sig
dess
benägna
förord
till
Kgl.
Majt
.
,
att
förberörda
regementsmöte
måtte
för
i
år
få
i
nåder
inställas
.

Sexmännen
visste
icke
närmare
någon
,
som
utan
församlingens
tillstånd
emottagit
inhysesfolk
från
andra
socknar
,
ävensom
de
ej
funnit
utsocknes
fattiga
besvära
socknen
med
tiggande
.
§
10
.

Modern
varnades
,
att
om
Gud
behagar
vidare
välsigna
henne
med
livsfrukt
,
hon
då
för
all
ting
må
akta
sig
för
vårdslöshet
om
sitt
foster
,
samt
tillsades
,
att
nästa
Söndag
sätta
sig
bak
i
kyrkan
,
då
hon
med
den
i
handboken
föreskrivna
bönen
från
Predikstolen
intages
till
församlingens
gemenskap
.
-
Så
vara
hänt
och
berättat
intyga
på
församlingens
vägnar
Carl
Fr
.

Maij
blev
allmän
Vallborgsm
.
Sockenstämma
hållen
med
St.
Malms
resp
.
församling
.
§
1
.

Prosten
sporde
vidare
,
om
icke
husmannen
Eric
Carlsson
i
Remrö
vore
därtill
skicklig
,
men
sockenmännen
svarade
,
att
denne
Eric
C
.
vore
mycket
sjuklig
,
bodde
nu
icke
i
Remrö
,
utan
i
Staksund
och
vore
således
långt
från
landsvägarna
,
samt
hade
ingen
hug
härför
.

Och
om
plåtbeslagens
anstrykande
lovade
Klockaren
Nylin
att
draga
försorg
.

Församlingen
hade
väl
kommit
överens
med
Eric
i
Remna
soldattorp
om
12
s
för
dagen
för
rödfärgningen
på
kyrkotaket
i
sommars
,
men
som
födan
var
dyr
och
han
farit
illa
med
sina
kläder
vid
detta
arbetet
,
så
beviljades
honom
dessutom
såsom
en
gåva
1
Rdr
32
s
.

Som
prosten
ofta
förnummit
,
att
en
stor
del
av
församlingens
ledamöter
tyckas
förglömt
,
vad
som
förr
beslutat
blivit
,
nämligen
att
ingen
har
lov
sitta
kvar
i
sockenstugan
eller
driva
på
Kyrkobacken
,
sedan
sammanringningen
skett
och
gudstjänsten
är
begynt
,
samt
ej
gå
ur
Kyrkan
,
förrän
allt
är
slutat
med
välsignelsen
;
så
upplästes
härom
§§
22
och
23
i
1784
års
protokoll
,
och
skulle
samma
§§
nästa
Bönedag
till
allas
underrättelse
å
predikstolen
uppläsas
.

In
fidem
protocolli
C
.
F
.
Maneck
Föregående
4
protokoll
är
upplästa
och
erkända
:

Sockenmännen
intygade
enhälligt
,
att
Brofogden
bättre
i
vår
,
än
förr
,
gjort
sin
syssla
,
så
att
inga
särdeles
svinpåtor
fanns
vid
Landsvägs
renarna
.
§
7
.

Skulle
åter
sammanskottet
ej
hinna
till
,
så
kommer
bristen
,
att
av
fattigkassan
fyllas
.

Resp
.
församlingen
kunde
ej
bifalla
,
att
Jan
Månssons
syster
i
Remna
,
en
änka
,
får
inflytta
i
socknen
.
§
11
.

Dessa
42
personer
fick
tillsammans
19
Rdr
24
sr
.
§
13
.

Sockenskräddare
ingav
skriftligen
sina
tankar
,
att
församlingen
borde
avskaffa
en
hop
överflödiga
modeller
på
kläder
ibland
allmogen
,
så
lydande
:
"
Som
här
uti
församlingen
är
ett
stort
överflöd
med
yppighet
uti
klädmodeller
,
och
som
nyfikenhet
av
skräddare
är
nog
orsaken
därtill
uti
början
;
alltså
har
socknens
hantverkare
kommit
överens
om
en
del
utav
dessa
modellers
borttagande
,
om
församlingens
hedervärda
allmoge
finner
sig
benägna
därtill
,
som
är
följande
.

Men
som
här
ännu
är
flera
,
som
icke
böra
tillåtas
,
att
intränga
sig
i
vår
profession
,
som
är
Eric
uti
Davidstorp
,
Pehr
i
Foglönäs
,
någon
Pehr
i
Ändebolshagstugan
och
son
Pehr
i
Byggslätten
,
samt
flera
utsocknes
intagande
,
och
som
detta
är
emot
Kungl.
författningar
,
hoppas
man
,
at
församlingen
ville
vara
så
goda
och
taga
det
i
övervägande
,
och
att
härefter
förekomma
flera
jämte
skräddare
,
har
vi
kommit
överens
,
att
ingen
skräddare
får
ha
någon
dräng
skriven
hos
sig
,
som
icke
är
i
hans
tjänst
,
vid
samma
vite
som
föresagt
är
.

Men
som
församlingen
befarade
,
att
summan
för
sådana
läkemedel
kunde
bli
nog
stor
för
kassan
att
bestrida
,
och
sade
sig
ej
heller
ha
råd
,
till
att
ytterligare
göra
pgr
sammanstkott
till
kassan
;
så
besvarades
frågan
med
nej
.

Sexmännen
anmodades
,
att
när
något
tjänstehjon
eller
inhyses
hjon
,
efter
hållet
husförhör
,
flyttar
till
annat
ställe
innom
socknen
,
ge
det
tillkänna
,
på
det
att
en
sådan
person
måtte
antecknas
i
husförhörsboken
vid
det
hemman
,
där
den
verkl
.
vistas
.
§
18
.

Dec
.
blev
allmän
Sockenstämma
hållen
med
St.
Malms
församlingen
,
då
följande
ärende
före
hades
:

De
beslöt
,
att
uppköpa
3
tolfter
plank
därtill
och
skulle
kyrkkassan
gå
i
förskott
för
betalningar
tills
vidare
.
§
11
.

Brofogden
hade
ingen
att
angiva
för
oringade
svinkreatur
§
3
.

In
fidem
C
.
F
.
Maneck
Föregående
2ne
protokoll
upplästes
i
allmän
Sockenstämma
d
.
6
.

Men
som
Klingström
nu
icke
var
närvarande
,
så
avgjordes
,
att
han
skulle
tillsägas
infinna
sig
i
sockenstug
.
nästa
Söndag
,
för
att
höras
häröver
.
§
6
.

Brofogden
uppgavs
ha
sitt
kall
väl
fullgjort
i
vår
och
anmodades
att
därmed
fortfara
.
§
4
.

I
anledning
av
1779
års
sockenstämmo
beslut
,
att
den
bonde
eller
torpare
,
som
till
Mickelsmässodanskalas
hållande
lämnar
sin
stuga
åt
tjänstefolk
och
annan
ungdom
,
skall
böta
3
Rdr
,
förklarade
sockenmännen
på
efterfrågan
,
det
meningen
då
varit
och
ännu
är
,
att
ej
heller
någon
soldat
på
sitt
torp
ägde
lämna
sin
stuga
eller
hus
till
ett
sådant
danskalas
,
utan
att
bli
till
ovannämnda
böter
förfallen
,
helst
mera
nämnda
beslut
eljest
skulle
bli
utan
allt
ändamål
,
och
soldaterna
ej
mer
än
andra
kunde
vara
berättigade
till
ordningars
befrämjande
och
underhållande
innom
församlingen
,
samt
att
orden
bonde
och
torpare
härvid
blivit
nyttjade
i
den
vidsträcktare
bemärkelse
,
vari
de
ofta
förekomma
,
det
förra
att
utmärka
innehavare
av
hemman
och
det
senare
åboer
å
oskattlagda
lägenheter
,
utan
avseende
för
övrigt
till
stånd
eller
näring
.
§
8
.

På
efterfrågan
sade
sexmännen
sig
icke
ha
hört
omtalas
,
att
något
Michelsm
.
danskalas
på
något
ställe
blivit
hållet
.

Torven
kunde
tagas
i
Prästgårdens
hagar
,
om
så
mycken
torv
täkt
där
finnes
.

Som
torv
tak
icke
länge
ha
bestånd
;
så
anhöll
Prosten
,
att
sockenmännen
täcktes
bestå
och
framdeles
på
torvtaken
över
bodar
och
brygghus
i
Prästgården
lägga
tegeltak
för
längre
varaktighet
skull
.

Prosten
,
som
förut
kände
församlingens
Herr
Patroni
gunstiga
bifall
till
nämnda
tegeltaks
påläggande
,
frågade
Befallningsman
Blomberg
vid
Djula
,
om
han
,
å
sitt
herrskaps
vägnar
,
samtyckte
till
hela
detta
sockenmännens
beslut
?

