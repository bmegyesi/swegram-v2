{"andra|NUM": "1", "arton|NUM": "1", "bakre|ADJ": "1", "brunch|NOUN": "1", "decimeter|NOUN": "1", "elva|NUM": "1", "ett|NUM": "1", "Europa|PROPN": "1", "fem|NUM": "1", "femte|NUM": "1", "femtio|NUM": "1", "femton|NUM": "1", "fjorton|NUM": "1", "fjärde|NUM": "1", "främre|ADJ": "1", "fyra|NUM": "1", "fyrtio|NUM": "1", "första|NUM": "1", "Grekland|PROPN": "1", "Göteborg|PROPN": "1", "hekto|NOUN": "1", "hela|NOUN": "1", "hundra|NUM": "1", "hundratusen|NUM": "1", "hörsel|NOUN": "1", "inrikesminister|NOUN": "1", "inrikespolitik|NOUN": "1", "Italien|PROPN": "1", "Kina|PROPN": "1", "kvällsmål|NOUN": "1", "känsel|NOUN": "1", "mellanmål|NOUN": "1", "miljard|NUM": "1", "miljon|NUM": "1", "milligram|NOUN": "1", "millimeter|NOUN": "1", "morbror|NOUN": "1", "månadsskifte|NOUN": "1", "nia|NOUN": "1", "nio|NUM": "1", "nionde|NUM": "1", "nittio|NUM": "1", "nitton|NUM": "1", "nordost|NOUN": "1", "Norge|PROPN": "1", "pingst|NOUN": "1", "Polen|PROPN": "1", "Ryssland|PROPN": "1", "sex|NUM": "1", "sexa|NOUN": "1", "sextio|NUM": "1", "sexton|NUM": "1", "sju|NUM": "1", "sjua|NOUN": "1", "sjunde|NUM": "1", "sjuttio|NUM": "1", "sjutton|NUM": "1", "sjätte|NUM": "1", "Stockholm|PROPN": "1", "storasyster|NOUN": "1", "Storbritannien|PROPN": "1", "syd|NOUN": "1", "sydväst|NOUN": "1", "sydöst|NOUN": "1", "syssling|NOUN": "1", "tia|NOUN": "1", "tio|NUM": "1", "tionde|NUM": "1", "tiotusen|NUM": "1", "tjugo|NUM": "1", "tolv|NUM": "1", "tre|NUM": "1", "tredje|NUM": "1", "trettio|NUM": "1", "tretton|NUM": "1", "tusen|NUM": "1", "två|NUM": "1", "utbildningsminister|NOUN": "1", "veckodag|NOUN": "1", "åtta|NOUN": "1", "åtta|NUM": "1", "åttio|NUM": "1", "åttonde|NUM": "1", "änkeman|NOUN": "1", "änkling|NOUN": "1", "ögonlock|NOUN": "1", "och (vardagl. å; förk. o.)|CCONJ": "1", "vara (vardagl. va)|VERB": "1", "i|ADP": "1", "ha|VERB": "1", "dess|PRON": "1", "det|PRON": "1", "en|DET": "1", "som|PRON": "1", "på|ADP": "1", "å|ADP": "1", "av|ADP": "1", "för|ADP": "1", "att|SCONJ": "1", "kunna|VERB": "1", "skola|AUX": "1", "jag|PRON": "1", "inte (formellt: icke, ej)|ADV": "1", "med|ADP": "1", "till|ADP": "1", "liten|ADJ": "1", "den|DET": "1", "ett|DET": "1", "analog|ADJ": "1", "unna|VERB": "1", "om|ADP": "1", "vi|PRON": "1", "men|CCONJ": "1", "man|PRON": "1", "de (vardagl. dom)|DET": "1", "få|VERB": "1", "så|ADV": "1", "som|CCONJ": "1", "sig (vardagl. sej)|PRON": "1", "han|PRON": "1", "de (vardagl. dom)|PRON": "1", "bli|VERB": "1", "komma|VERB": "1", "det|DET": "1", "sin|PRON": "1", "eller|CCONJ": "1", "från|ADP": "1", "mycket|ADV": "1", "vilja|VERB": "1", "all|PRON": "1", "göra|VERB": "1", "om|SCONJ": "1", "annan|PRON": "1", "du|PRON": "1", "någon (vardagl. nån, förk. ngn)|PRON": "1", "finna|VERB": "1", "ta (el. taga)|VERB": "1", "när|ADV": "1", "se|VERB": "1", "måste|AUX": "1", "detta|PRON": "1", "stor|ADJ": "1", "nu|ADV": "1", "gå|VERB": "1", "säga|VERB": "1", "den|PRON": "1", "vad (vardagl. va)|PRON": "1", "år|NOUN": "1", "äga|VERB": "1", "under|ADP": "1", "betyda|VERB": "1", "också (vardagl. oxå)|ADV": "1", "där|ADV": "1", "då|ADV": "1", "min|PRON": "1", "böra|AUX": "1", "hur|ADV": "1", "mig (vardagl. mej)|PRON": "1", "mot|ADP": "1", "bara|ADV": "1", "vilken|PRON": "1", "ut|ADV": "1", "ny|ADJ": "1", "vid|ADP": "1", "än|CCONJ": "1", "bra|ADJ": "1", "ingen|PRON": "1", "dem (vardagl. dom)|PRON": "1", "efter|ADP": "1", "upp|PART": "1", "hon|PRON": "1", "lite|ADV": "1", "denna|PRON": "1", "in|ADV": "1", "mycket|ADJ": "1", "över|ADP": "1", "ge (formellt giva)|VERB": "1", "vår (vardagl. våran)|PRON": "1", "del|NOUN": "1", "här|ADV": "1", "även|ADV": "1", "skriva|VERB": "1", "tid|NOUN": "1", "ju|ADV": "1", "sedan (vardagl. sen)|ADV": "1", "te sig|VERB": "1", "riva|VERB": "1", "börja|VERB": "1", "hel|ADJ": "1", "dag|NOUN": "1", "själv|PRON": "1", "människa|NOUN": "1", "land|NOUN": "1", "svensk|ADJ": "1", "fråga|NOUN": "1", "oss|PRON": "1", "tro|VERB": "1", "el|NOUN": "1", "tycka|VERB": "1", "kommentar|NOUN": "1", "veta|VERB": "1", "idag (el. i dag)|ADV": "1", "försöka|VERB": "1", "behöva|VERB": "1", "samma|PRON": "1", "mellan|ADP": "1", "känna|VERB": "1", "läsa|VERB": "1", "ro|VERB": "1", "kanske|ADV": "1", "lik|ADJ": "1", "låta|VERB": "1", "olik|ADJ": "1", "sådan|PRON": "1", "sätt|NOUN": "1", "hans|PRON": "1", "din|PRON": "1", "gång|NOUN": "1", "stå|VERB": "1", "inom|ADP": "1", "visa|VERB": "1", "använda|VERB": "1", "vända|VERB": "1", "hålla|VERB": "1", "genom|ADP": "1", "helt|ADV": "1", "fler|ADJ": "1", "utan|ADP": "1", "väl|ADV": "1", "barn|NOUN": "1", "enligt|ADP": "1", "tänka|VERB": "1", "ni|PRON": "1", "viktig|ADJ": "1", "ring|NOUN": "1", "eftersom|SCONJ": "1", "liv|NOUN": "1", "deras|PRON": "1", "värld|NOUN": "1", "viss|ADJ": "1", "dock|ADV": "1", "egen|ADJ": "1", "folk|NOUN": "1", "regering|NOUN": "1", "fram|PART": "1", "honom|PRON": "1", "söka|VERB": "1", "dig (vardagl. dej)|PRON": "1", "utan|CCONJ": "1", "sak|NOUN": "1", "hög|ADJ": "1", "länge|ADV": "1", "person|NOUN": "1", "ligga|VERB": "1", "son|NOUN": "1", "både|CCONJ": "1", "just|ADV": "1", "lägga|VERB": "1", "antal|NOUN": "1", "redan|ADV": "1", "kvinna|NOUN": "1", "problem|NOUN": "1", "fall|NOUN": "1", "man|NOUN": "1", "aldrig|ADV": "1", "ofta|ADV": "1", "varje|DET": "1", "artikel|NOUN": "1", "anse|VERB": "1", "öva|VERB": "1", "lag|NOUN": "1", "slag|NOUN": "1", "tal|NOUN": "1", "åt|ADP": "1", "nog|ADV": "1", "bok|NOUN": "1", "varför|ADV": "1", "handla|VERB": "1", "gammal|ADJ": "1", "bild|NOUN": "1", "sida|NOUN": "1", "så|SCONJ": "1", "öka|VERB": "1", "därför|ADV": "1", "sen|ADJ": "1", "god|ADJ": "1", "hos|ADP": "1", "alltid|ADV": "1", "skapa|VERB": "1", "arbete|NOUN": "1", "kapa|VERB": "1", "samt|CCONJ": "1", "blogg|NOUN": "1", "innan|SCONJ": "1", "som|ADV": "1", "ur|ADP": "1", "gälla|VERB": "1", "verka|VERB": "1", "tala|VERB": "1", "bära|VERB": "1", "för|ADV": "1", "väg|NOUN": "1", "samhälle|NOUN": "1", "alltså|ADV": "1", "stat|NOUN": "1", "stad|NOUN": "1", "höra|VERB": "1", "innebära|VERB": "1", "genom att|SCONJ": "1", "företag|NOUN": "1", "möjlighet|NOUN": "1", "ord|NOUN": "1", "politisk|ADJ": "1", "välja|VERB": "1", "er|PRON": "1", "förstå|VERB": "1", "inlägg|NOUN": "1", "ägg|NOUN": "1", "te|NOUN": "1", "spela|VERB": "1", "så att|SCONJ": "1", "lika|ADV": "1", "hitta|VERB": "1", "tag|NOUN": "1", "dra|VERB": "1", "leda|VERB": "1", "gärna|ADV": "1", "ändå|ADV": "1", "förslag|NOUN": "1", "lyckas|VERB": "1", "dessutom|ADV": "1", "område|NOUN": "1", "svår|ADJ": "1", "lära|VERB": "1", "sätta|VERB": "1", "plats|NOUN": "1", "lång|ADJ": "1", "lämna|VERB": "1", "bygga|VERB": "1", "politik|NOUN": "1", "tidigare|ADV": "1", "kalla|VERB": "1", "peng|NOUN": "1", "väldigt|ADV": "1", "leva|VERB": "1", "ställa|VERB": "1", "följa|VERB": "1", "vecka|NOUN": "1", "ja|INTJ": "1", "ske|VERB": "1", "parti|NOUN": "1", "kräva|VERB": "1", "utveckling|NOUN": "1", "faktiskt|ADV": "1", "ena|VERB": "1", "svara|VERB": "1", "ner|PART": "1", "fortsätta|VERB": "1", "skola|NOUN": "1", "bruka|VERB": "1", "mål|NOUN": "1", "par|NOUN": "1", "sent|ADV": "1", "ekonomisk|ADJ": "1", "kl. (klockan)|NOUN": "1", "dålig|ADJ": "1", "namn|NOUN": "1", "igen|ADV": "1", "verkligen|ADV": "1", "mena|VERB": "1", "fortfarande|ADV": "1", "grupp|NOUN": "1", "beslut|NOUN": "1", "även om|SCONJ": "1", "enda|ADJ": "1", "bort|PART": "1", "slå|VERB": "1", "möjlig|ADJ": "1", "många|PRON": "1", "hända|VERB": "1", "ämna|AUX": "1", "endast|ADV": "1", "miljon|NOUN": "1", "vidare|ADV": "1", "ganska|ADV": "1", "svar|NOUN": "1", "varenda|DET": "1", "istället (el. i stället)|ADV": "1", "först|ADV": "1", "arbeta|VERB": "1", "heller|ADV": "1", "riktigt|ADV": "1", "hand|NOUN": "1", "uppgift|NOUN": "1", "fungera (vardagl. funka)|VERB": "1", "beta|VERB": "1", "köpa|VERB": "1", "nästan|ADV": "1", "bra|ADV": "1", "bland|ADP": "1", "december|NOUN": "1", "sitta|VERB": "1", "precis|ADV": "1", "hennes|PRON": "1", "åta sig|VERB": "1", "bland annat (förk. bl.a.)|ADV": "1", "krig|NOUN": "1", "till exempel (förk. t.ex., t ex)|ADV": "1", "tillsammans|ADV": "1", "henne|PRON": "1", "intressant|ADJ": "1", "val|NOUN": "3", "kyrka|NOUN": "1", "egentligen|ADV": "1", "inför|ADP": "1", "historia|NOUN": "1", "jobb|NOUN": "1", "berätta|VERB": "1", "vanlig|ADJ": "1", "rätta|VERB": "1", "januari|NOUN": "1", "information|NOUN": "1", "flest|ADJ": "1", "ung|ADJ": "1", "en|PRON": "1", "tillbaka (vardagl. tillbaks)|PART": "1", "film|NOUN": "1", "ibland (el. i bland)|ADV": "1", "medan (vardagl. medans)|SCONJ": "1", "slut|NOUN": "1", "massa|NOUN": "1", "tanke|NOUN": "1", "akt|NOUN": "1", "procent|NOUN": "1", "månad|NOUN": "1", "sista|ADJ": "1", "ätt|NOUN": "1", "sluta|VERB": "1", "verksamhet|NOUN": "1", "rätt|NOUN": "1", "samtidigt|ADV": "1", "emot|ADP": "1", "stöd|NOUN": "1", "familj|NOUN": "1", "vem|PRON": "1", "åka|VERB": "1", "betala|VERB": "1", "kommun|NOUN": "1", "resultat|NOUN": "1", "utveckla|VERB": "1", "föra|VERB": "1", "hjälpa|VERB": "1", "nästa|ADJ": "1", "nära|ADV": "1", "nej|INTJ": "1", "text|NOUN": "1", "exempel|NOUN": "1", "särskilt|ADV": "1", "debatt|NOUN": "1", "när det gäller|ADP": "1", "på grund av (förk. p.g.a, pga., p g a)|ADV": "1", "situation|NOUN": "1", "europeisk|ADJ": "1", "form|NOUN": "1", "orm|NOUN": "1", "råd|NOUN": "1", "november|NOUN": "1", "makt|NOUN": "1", "social|ADJ": "1", "vinna|VERB": "1", "kvar|PART": "1", "system|NOUN": "1", "vänta|VERB": "1", "tidig|ADJ": "1", "åtgärd|NOUN": "1", "krav|NOUN": "1", "skillnad|NOUN": "1", "riksdag|NOUN": "1", "internationell|ADJ": "1", "nationell|ADJ": "1", "jobba|VERB": "1", "klara|VERB": "1", "typ|NOUN": "1", "kring|ADP": "1", "båda (vardagl. bägge)|PRON": "1", "cirka (förk. ca)|ADV": "1", "tur|NOUN": "1", "polis|NOUN": "1", "medium|NOUN": "1", "låg|ADJ": "1", "varandra (vardagl. varann)|PRON": "1", "mun|NOUN": "1", "ansvar|NOUN": "1", "roll|NOUN": "1", "regel|NOUN": "1", "oktober|NOUN": "1", "prata|VERB": "1", "organisation|NOUN": "1", "medlem|NOUN": "1", "fråga|VERB": "1", "anmäla|VERB": "1", "nå|VERB": "1", "bo|VERB": "1", "krona|NOUN": "1", "stämma|VERB": "1", "rättighet|NOUN": "1", "sedan (vardagl. sen)|ADP": "1", "bakom|ADP": "1", "efter att|SCONJ": "1", "därmed|ADV": "1", "med|ADV": "1", "hus|NOUN": "1", "vän|NOUN": "1", "dela|VERB": "1", "februari|NOUN": "1", "kort|ADJ": "1", "grund|NOUN": "1", "runt|ADP": "1", "framtid|NOUN": "1", "köra|VERB": "1", "etikett|NOUN": "1", "fri|ADJ": "1", "behov|NOUN": "1", "timme (el. timma)|NOUN": "1", "september|NOUN": "1", "hoppas|VERB": "1", "ensam|ADJ": "1", "snart|ADV": "1", "rätt|ADV": "1", "förklara|VERB": "1", "ledning|NOUN": "1", "intresse|NOUN": "1", "tvinga|VERB": "1", "påverka|VERB": "1", "anledning|NOUN": "1", "titta|VERB": "1", "minska|VERB": "1", "i alla fall (el. iallafall; förk. iaf)|ADV": "1", "däremot|ADV": "1", "direkt|ADV": "1", "ekonomi|NOUN": "1", "bestämma|VERB": "1", "skicka|VERB": "1", "trots|ADP": "1", "åsikt|NOUN": "1", "diskussion|NOUN": "1", "rad|NOUN": "1", "faktum|NOUN": "1", "tidning|NOUN": "1", "mening|NOUN": "1", "utanför|ADP": "1", "rätt|ADJ": "1", "gemensam|ADJ": "1", "klar|ADJ": "1", "juni|NOUN": "1", "is|NOUN": "1", "bil|NOUN": "1", "myndighet|NOUN": "1", "nummer (förk. nr)|NOUN": "1", "allmän|ADJ": "1", "musik|NOUN": "1", "ändra|VERB": "1", "träffa|VERB": "1", "ihop|PART": "1", "diskutera|VERB": "1", "driva|VERB": "1", "sälja|VERB": "1", "sakna|VERB": "1", "program|NOUN": "1", "ifrån|ADP": "1", "länka|VERB": "1", "kunskap|NOUN": "1", "snabbt|ADV": "1", "maj|NOUN": "1", "amerikansk|ADJ": "1", "tyda|VERB": "1", "särskild|ADJ": "1", "början|NOUN": "1", "naturligtvis|ADV": "1", "skäl|NOUN": "1", "fin|ADJ": "1", "genomföra|VERB": "1", "liksom|ADV": "1", "via|ADP": "1", "före|ADP": "1", "dom|NOUN": "1", "risk|NOUN": "1", "enkel|ADJ": "1", "alls|ADV": "1", "pris|NOUN": "1", "räkna|VERB": "1", "beskriva|VERB": "1", "hem|PART": "1", "möta|VERB": "1", "såsom|SCONJ": "1", "idé|NOUN": "1", "gram|NOUN": "1", "förra|ADJ": "1", "tjänst|NOUN": "1", "heta|VERB": "1", "kultur|NOUN": "1", "äta|VERB": "1", "syfte|NOUN": "1", "princip|NOUN": "1", "flytta|VERB": "1", "ute|ADV": "1", "utgöra|VERB": "1", "politiker|NOUN": "1", "lätt|ADJ": "1", "förälder|NOUN": "1", "marknad|NOUN": "1", "nämligen|ADV": "1", "tydlig|ADJ": "1", "utbildning|NOUN": "1", "röra|VERB": "1", "nivå|NOUN": "1", "april|NOUN": "1", "mängd|NOUN": "1", "betydelse|NOUN": "1", "kristen|ADJ": "1", "dö|VERB": "1", "mars|NOUN": "1", "allt|ADV": "1", "kväll|NOUN": "1", "bildning|NOUN": "1", "länk|NOUN": "1", "växa|VERB": "1", "per|ADP": "1", "offentlig|ADJ": "1", "såväl|CCONJ": "1", "våga|VERB": "1", "vatten|NOUN": "1", "håll|NOUN": "1", "mänsklig|ADJ": "1", "demokrati|NOUN": "1", "fatta|VERB": "1", "jord|NOUN": "1", "känsla|NOUN": "1", "förändring|NOUN": "1", "nämna|VERB": "1", "tyvärr|ADV": "1", "enskild|ADJ": "1", "rätt|PART": "1", "be (el. bedja)|VERB": "1", "punkt|NOUN": "1", "ändring|NOUN": "1", "mission|NOUN": "1", "igår (el. i går)|ADV": "1", "kommission|NOUN": "1", "ort|NOUN": "1", "anta|VERB": "1", "trots att|SCONJ": "1", "spel|NOUN": "1", "språk|NOUN": "1", "föreslå|VERB": "1", "igenom|ADP": "1", "undra|VERB": "1", "eget|ADJ": "1", "möte|NOUN": "1", "mat|NOUN": "1", "gräns|NOUN": "1", "lyssna|VERB": "1", "delta|VERB": "1", "samarbete|NOUN": "1", "annars|ADV": "1", "falla|VERB": "1", "nära|ADJ": "1", "rum|NOUN": "1", "ungefär|ADV": "1", "starta|VERB": "1", "inse|VERB": "1", "internet|NOUN": "1", "hov|NOUN": "1", "öppen|ADJ": "1", "bidra|VERB": "1", "död|NOUN": "1", "luta|VERB": "1", "öga|NOUN": "1", "säkert|ADV": "1", "ämne|NOUN": "1", "få|ADJ": "1", "augusti|NOUN": "1", "socialdemokrat (vardagl. sosse)|NOUN": "1", "projekt|NOUN": "1", "övrig|ADJ": "1", "dels|CCONJ": "1", "framför allt (el. framförallt)|ADV": "1", "positiv|ADJ": "1", "rolig|ADJ": "1", "port|NOUN": "1", "bero|VERB": "1", "kropp|NOUN": "1", "minnas|VERB": "1", "handling|NOUN": "1", "rösta|VERB": "1", "riktig|ADJ": "1", "rapport|NOUN": "1", "lösning|NOUN": "1", "personlig|ADJ": "1", "kommentera|VERB": "1", "som att|SCONJ": "1", "gilla|VERB": "1", "bryta|VERB": "1", "hjälp|NOUN": "1", "juli|NOUN": "1", "innehålla|VERB": "1", "liknande|ADJ": "1", "tillfälle|NOUN": "1", "inte ens|ADV": "1", "känd|ADJ": "1", "forskning|NOUN": "1", "kraft|NOUN": "1", "helt enkelt|ADV": "1", "brott|NOUN": "1", "exempelvis|ADV": "1", "röst|NOUN": "1", "bjuda|VERB": "1", "till och med (förk. t.o.m., t o m)|ADV": "1", "hävda|VERB": "1", "hamna|VERB": "1", "effekt|NOUN": "1", "enhet|NOUN": "1", "det vill säga (förk. d.v.s., dvs.)|ADV": "1", "kontakt|NOUN": "1", "takt|NOUN": "1", "värde|NOUN": "1", "förutsättning|NOUN": "1", "sats|NOUN": "1", "medlemsstat|NOUN": "1", "hinna|VERB": "1", "sanning|NOUN": "1", "religion|NOUN": "1", "källa|NOUN": "1", "må|VERB": "1", "kostnad|NOUN": "1", "medborgare|NOUN": "1", "förhållande|NOUN": "1", "far (el. fader, vardagl. farsa)|NOUN": "1", "miljard|NOUN": "1", "ungdom|NOUN": "1", "släppa|VERB": "1", "enbart|ADV": "1", "drag|NOUN": "1", "verklighet|NOUN": "1", "författare|NOUN": "1", "tillgång|NOUN": "1", "nödvändig|ADJ": "1", "full|ADJ": "1", "frihet|NOUN": "1", "passa|VERB": "1", "lokal|ADJ": "1", "ytterligare|ADV": "1", "öppna|VERB": "1", "införa|VERB": "1", "ledare|NOUN": "1", "mamma|NOUN": "1", "sammanhang|NOUN": "1", "svensk|NOUN": "1", "hemma|ADV": "1", "produkt|NOUN": "1", "därefter|ADV": "1", "efter|ADV": "1", "match|NOUN": "1", "tro|NOUN": "1", "alldeles|ADV": "1", "lätt|ADV": "1", "sann|ADJ": "1", "uppfattning|NOUN": "1", "demokrat|NOUN": "1", "bolag|NOUN": "1", "erfarenhet|NOUN": "1", "kritik|NOUN": "1", "grad|NOUN": "1", "jude|NOUN": "1", "vacker|ADJ": "1", "erbjuda|VERB": "1", "kamp|NOUN": "1", "period|NOUN": "1", "modern|ADJ": "1", "spelare|NOUN": "1", "elev|NOUN": "1", "utredning|NOUN": "1", "ingå|VERB": "1", "kung|NOUN": "1", "bestå|VERB": "1", "katt|NOUN": "1", "konstatera|VERB": "1", "dit|ADV": "1", "klart|ADV": "1", "nuvarande|ADJ": "1", "styra|VERB": "1", "förlora|VERB": "1", "vit|ADJ": "1", "klocka|NOUN": "1", "påstå|VERB": "1", "skatt|NOUN": "1", "besluta|VERB": "1", "befolkning|NOUN": "1", "avse|VERB": "1", "ro|NOUN": "1", "privat|ADJ": "1", "steg|NOUN": "1", "art|NOUN": "1", "stödja|VERB": "1", "ond|ADJ": "1", "plan|NOUN": "2", "resa|NOUN": "1", "utom|ADP": "1", "hund|NOUN": "1", "syn|NOUN": "1", "glömma|VERB": "1", "avtal|NOUN": "1", "lek|NOUN": "1", "kul|ADJ": "1", "natt|NOUN": "1", "förändra|VERB": "1", "ange|VERB": "1", "någonting|PRON": "1", "förstås|ADV": "1", "individ|NOUN": "1", "älska|VERB": "1", "motion|NOUN": "1", "glad|ADJ": "1", "ned|PART": "1", "dator|NOUN": "1", "miljö|NOUN": "1", "ek|NOUN": "1", "åtminstone|ADV": "1", "presentera|VERB": "1", "stanna|VERB": "1", "byta|VERB": "1", "alternativ|NOUN": "1", "minut|NOUN": "1", "ingenting|PRON": "1", "uppleva|VERB": "1", "samla|VERB": "1", "svart|ADJ": "1", "bakgrund|NOUN": "1", "skott|NOUN": "1", "ö|NOUN": "1", "kärlek|NOUN": "1", "metod|NOUN": "1", "äldre|ADJ": "1", "säker|ADJ": "1", "borgare|NOUN": "1", "gud|NOUN": "1", "insats|NOUN": "1", "tysk|ADJ": "1", "kontroll|NOUN": "1", "lösa|VERB": "1", "kolla|VERB": "1", "fylla|VERB": "1", "bestämmelse|NOUN": "1", "ris|NOUN": "1", "drabba|VERB": "1", "nät|NOUN": "1", "teknik|NOUN": "1", "resurs|NOUN": "1", "försök|NOUN": "1", "fara|VERB": "1", "tjäna|VERB": "1", "argument|NOUN": "1", "behandla|VERB": "1", "ren|ADJ": "1", "fru|NOUN": "1", "sjuk|ADJ": "1", "istället för (el. i stället för)|ADP": "1", "våld|NOUN": "1", "utföra|VERB": "1", "ställning|NOUN": "1", "främst|ADV": "1", "räcka|VERB": "1", "bättre|ADV": "1", "fundera|VERB": "1", "visst|ADV": "1", "sommar|NOUN": "1", "rörelse|NOUN": "1", "kund|NOUN": "1", "villkor|NOUN": "1", "tillbaka (vardagl. tillbaks)|ADV": "1", "högt|ADV": "1", "president|NOUN": "1", "emellertid|ADV": "1", "händelse|NOUN": "1", "uppstå|VERB": "1", "acceptera|VERB": "1", "huvud|NOUN": "1", "sök|NOUN": "1", "snabb|ADJ": "1", "så kallad (förk. s.k., s k)|ADV": "1", "framför|ADP": "1", "ande|NOUN": "1", "bilda|VERB": "1", "orsak|NOUN": "1", "försvinna|VERB": "1", "fel|NOUN": "1", "innehåll|NOUN": "1", "natur|NOUN": "1", "begrepp|NOUN": "1", "för att|SCONJ": "1", "konflikt|NOUN": "1", "tack|INTJ": "1", "djur|NOUN": "1", "chans|NOUN": "1", "samtidigt som|SCONJ": "1", "demokratisk|ADJ": "1", "fel|ADV": "1", "läge|NOUN": "1", "sprida|VERB": "1", "växt|NOUN": "1", "förutom|ADP": "1", "i samband med|ADP": "1", "styck|NOUN": "1", "utskott|NOUN": "1", "muslim|NOUN": "1", "ordning|NOUN": "1", "uppdrag|NOUN": "1", "mark|NOUN": "1", "säkerhet|NOUN": "1", "linje|NOUN": "1", "bank|NOUN": "1", "önska|VERB": "1", "givetvis|ADV": "1", "studie|NOUN": "1", "fredag|NOUN": "1", "lärare|NOUN": "1", "statlig|ADJ": "1", "söndag|NOUN": "1", "fel|ADJ": "1", "speciellt|ADV": "1", "röd|ADJ": "1", "television (el. teve, tv)|NOUN": "1", "hot|NOUN": "1", "verk|NOUN": "1", "publicera|VERB": "1", "stund|NOUN": "1", "tillhöra|VERB": "1", "omfatta|VERB": "1", "material|NOUN": "1", "pelare|NOUN": "1", "hjärta|NOUN": "1", "knappast|ADV": "1", "befinna|VERB": "1", "part|NOUN": "1", "trevlig|ADJ": "1", "höst|NOUN": "1", "skilja|VERB": "1", "ens|ADV": "1", "förmåga|NOUN": "1", "döda|VERB": "1", "stånd|NOUN": "1", "peka|VERB": "1", "bedömning|NOUN": "1", "ringa|VERB": "1", "betrakta|VERB": "1", "by|NOUN": "1", "utifrån|ADP": "1", "brist|NOUN": "1", "hänga|VERB": "1", "tillräckligt|ADV": "1", "måndag|NOUN": "1", "aktuell|ADJ": "1", "någonsin (vardagl. nånsin)|ADV": "1", "tillåta|VERB": "1", "universitet|NOUN": "1", "konsekvens|NOUN": "1", "ställe|NOUN": "1", "hård|ADJ": "1", "majoritet|NOUN": "1", "domstol|NOUN": "1", "ordförande|NOUN": "1", "lördag|NOUN": "1", "låt|NOUN": "1", "herr|NOUN": "1", "sekvens|NOUN": "1", "förekomma|VERB": "1", "stoppa|VERB": "1", "nyhet|NOUN": "1", "journalist|NOUN": "1", "kris|NOUN": "1", "rycka|VERB": "1", "trycka|VERB": "1", "betydligt|ADV": "1", "kosta|VERB": "1", "band|NOUN": "1", "numera (el. numer)|ADV": "1", "tillstånd|NOUN": "1", "värd|ADJ": "1", "igen|PART": "1", "imorgon (el. i morgon)|ADV": "1", "klass|NOUN": "1", "uttrycka|VERB": "1", "slutsats|NOUN": "1", "global|ADJ": "1", "mitt|ADV": "1", "stol|NOUN": "1", "ytterligare|ADJ": "1", "effektiv|ADJ": "1", "resa|VERB": "1", "förbättra|VERB": "1", "rädda|VERB": "1", "list|NOUN": "1", "relation|NOUN": "1", "agera|VERB": "1", "central|ADJ": "1", "flera|PRON": "1", "undersökning|NOUN": "1", "uppnå|VERB": "1", "krona (förk. kr.)|NOUN": "1", "perspektiv|NOUN": "1", "plötsligt|ADV": "1", "naturlig|ADJ": "1", "ålder|NOUN": "1", "process|NOUN": "1", "uttryck|NOUN": "1", "lista|NOUN": "1", "allra|ADV": "1", "sökning|NOUN": "1", "ökning|NOUN": "1", "därför att|SCONJ": "1", "rysk|ADJ": "1", "jämföra (förk. jfr)|VERB": "1", "tills|SCONJ": "1", "intresserad|ADJ": "1", "totalt|ADV": "1", "hantera|VERB": "1", "förvänta|VERB": "1", "medel|NOUN": "1", "vika|VERB": "1", "döma|VERB": "1", "besöka|VERB": "1", "hem|NOUN": "1", "var|ADV": "1", "täcka|VERB": "1", "borgerlig|ADJ": "1", "inleda|VERB": "1", "helg|NOUN": "1", "undvika|VERB": "1", "ryck|NOUN": "1", "tryck|NOUN": "1", "tydligen|ADV": "1", "aktiv|ADJ": "1", "höja|VERB": "1", "pappa|NOUN": "1", "varkeneller|CCONJ": "1", "religiös|ADJ": "1", "råka|VERB": "1", "verklig|ADJ": "1", "rent|ADV": "1", "fantastisk|ADJ": "1", "grundläggande|ADJ": "1", "upptäcka|VERB": "1", "erkänna|VERB": "1", "helig|ADJ": "1", "lön|NOUN": "1", "historisk|ADJ": "1", "rest|NOUN": "1", "halv|ADJ": "1", "andel|NOUN": "1", "besök|NOUN": "1", "teknisk|ADJ": "1", "kasta|VERB": "1", "hemsida|NOUN": "1", "bedöma|VERB": "1", "torsdag|NOUN": "1", "tillväxt|NOUN": "1", "läsare|NOUN": "1", "forskare|NOUN": "1", "bidrag|NOUN": "1", "onsdag|NOUN": "1", "vilja|NOUN": "1", "sol|NOUN": "1", "inte minst|ADV": "1", "analys|NOUN": "1", "ovan|ADV": "1", "lagstiftning|NOUN": "1", "militär|ADJ": "1", "toppa|VERB": "1", "sort|NOUN": "1", "fördel|NOUN": "1", "skydda|VERB": "1", "nyttja|VERB": "1", "utnyttja|VERB": "1", "teori|NOUN": "1", "fransk|ADJ": "1", "pågå|VERB": "1", "samling|NOUN": "1", "flertal|NOUN": "1", "snarare|ADV": "1", "försvara|VERB": "1", "modell|NOUN": "1", "skön|ADJ": "1", "vapen|NOUN": "1", "således|ADV": "1", "förening|NOUN": "1", "lyfta|VERB": "1", "eftermiddag (förk. em.)|NOUN": "1", "soldat|NOUN": "1", "märka|VERB": "1", "gemenskap|NOUN": "1", "ösa|VERB": "1", "fast|CCONJ": "1", "styrka|NOUN": "1", "ersätta|VERB": "1", "kille|NOUN": "1", "vård|NOUN": "1", "fullt|ADV": "1", "ägna|VERB": "1", "oavsett|ADP": "1", "poäng|NOUN": "1", "satsa|VERB": "1", "moderat|NOUN": "1", "rida|VERB": "1", "jo|INTJ": "1", "tisdag|NOUN": "1", "död|ADJ": "1", "allmänt|ADV": "1", "avsluta|VERB": "1", "sova|VERB": "1", "inne|ADV": "1", "flicka|NOUN": "1", "sedan (vardagl. sen)|SCONJ": "1", "total|ADJ": "1", "allvarlig|ADJ": "1", "fram|ADV": "1", "ljus|NOUN": "1", "sjukdom|NOUN": "1", "unge|NOUN": "1", "i form av|ADP": "1", "vikt|NOUN": "1", "rik|ADJ": "1", "region|NOUN": "1", "samtal|NOUN": "1", "negativ|ADJ": "1", "mycket|PRON": "1", "i år|ADV": "1", "igång|PART": "1", "vändning|NOUN": "1", "antingeneller|CCONJ": "1", "föda|VERB": "1", "åter|ADV": "1", "arbetare|NOUN": "1", "skjuta|VERB": "1", "tradition|NOUN": "1", "hämta|VERB": "1", "församling|NOUN": "1", "hav|NOUN": "1", "energi|NOUN": "1", "bred|ADJ": "1", "vad gäller|ADP": "1", "fast|PART": "1", "påpeka|VERB": "1", "bättra|VERB": "1", "skaffa|VERB": "1", "utgå|VERB": "1", "samtlig|ADJ": "1", "stärka|VERB": "1", "läkare|NOUN": "1", "fattig|ADJ": "1", "grepp|NOUN": "1", "hej|INTJ": "1", "utsätta|VERB": "1", "spännande|ADJ": "1", "fort|ADV": "1", "sikt|NOUN": "1", "revolution|NOUN": "1", "brev|NOUN": "1", "personal|NOUN": "1", "skada|NOUN": "1", "illa|ADV": "1", "kämpa|VERB": "1", "alltför|ADV": "1", "tecken|NOUN": "1", "siffra|NOUN": "1", "tydligt|ADV": "1", "än (el. ännu)|ADV": "1", "hårt|ADV": "1", "absolut|ADV": "1", "eka|VERB": "1", "engelsk|ADJ": "1", "praktik|NOUN": "1", "förmodligen|ADV": "1", "hoppa|VERB": "1", "morgon|NOUN": "1", "tjej|NOUN": "1", "konstig|ADJ": "1", "union|NOUN": "1", "kommande|ADJ": "1", "avgöra|VERB": "1", "chef|NOUN": "1", "vis|NOUN": "1", "strid|NOUN": "1", "sända|VERB": "1", "missa|VERB": "1", "bedriva|VERB": "1", "etcetera (el. et cetera, förk. etc.)|ADV": "1", "anföra|VERB": "1", "varm|ADJ": "1", "hit|ADV": "1", "berättelse|NOUN": "1", "produktion|NOUN": "1", "kapitel (förk. kap.)|NOUN": "1", "hindra|VERB": "1", "konst|NOUN": "1", "speciell|ADJ": "1", "allvar|NOUN": "1", "grön|ADJ": "1", "vår|NOUN": "1", "meddela|VERB": "1", "omöjlig|ADJ": "1", "tillämpa|VERB": "1", "skydd|NOUN": "1", "hittills|ADV": "1", "sällan|ADV": "1", "position|NOUN": "1", "behandling|NOUN": "1", "omfattande|ADJ": "1", "skog|NOUN": "1", "kritisera|VERB": "1", "förklaring|NOUN": "1", "springa|VERB": "1", "oerhört|ADV": "1", "uppfatta|VERB": "1", "foto|NOUN": "1", "islam|NOUN": "1", "stänga|VERB": "1", "aning|NOUN": "1", "försvar|NOUN": "1", "meter|NOUN": "1", "evolution|NOUN": "1", "funktion|NOUN": "1", "dotter|NOUN": "1", "värdering|NOUN": "1", "råda|VERB": "1", "ersättning|NOUN": "1", "slippa|VERB": "1", "självklart|ADV": "1", "lämplig|ADJ": "1", "ting|NOUN": "1", "minne|NOUN": "1", "strategi|NOUN": "1", "dyka|VERB": "1", "orka|VERB": "1", "kontrollera|VERB": "1", "planera|VERB": "1", "färg|NOUN": "1", "lova|VERB": "1", "citera|VERB": "1", "finansiell|ADJ": "1", "ständigt|ADV": "1", "spår|NOUN": "1", "kall|ADJ": "1", "vuxen|ADJ": "1", "allians|NOUN": "1", "faktor|NOUN": "1", "kvalitet (el. kvalité)|NOUN": "1", "upp|ADV": "1", "utländsk|ADJ": "1", "svag|ADJ": "1", "sköta|VERB": "1", "vägra|VERB": "1", "rike|NOUN": "1", "framgå|VERB": "1", "judisk|ADJ": "1", "studera|VERB": "1", "farlig|ADJ": "1", "framgång|NOUN": "1", "tolka|VERB": "1", "billig|ADJ": "1", "iväg|PART": "1", "student|NOUN": "1", "och så vidare (förk. o.s.v., osv.)|ADV": "1", "visserligen|ADV": "1", "vara|NOUN": "1", "undantag|NOUN": "1", "tillgänglig|ADJ": "1", "enorm|ADJ": "1", "behålla|VERB": "1", "dricka|VERB": "1", "aktion|NOUN": "1", "bry sig|VERB": "1", "relativt|ADV": "1", "tung|ADJ": "1", "arbetsgivare|NOUN": "1", "med hjälp av|ADP": "1", "tvärtom (el. tvärt om)|ADV": "1", "notera|VERB": "1", "nation|NOUN": "1", "sänka|VERB": "1", "ärende|NOUN": "1", "givare|NOUN": "1", "kull|NOUN": "1", "nyligen|ADV": "1", "rättelse|NOUN": "1", "delvis|ADV": "1", "medföra|VERB": "1", "ifrågasätta|VERB": "1", "för övrigt|ADV": "1", "län|NOUN": "1", "gata|NOUN": "1", "medveten|ADJ": "1", "serie|NOUN": "1", "rimlig|ADJ": "1", "ty|CCONJ": "1", "invandrare|NOUN": "1", "dörr|NOUN": "1", "direktiv|NOUN": "1", "stiga|VERB": "1", "tiga|VERB": "1", "fot|NOUN": "1", "begränsad|ADJ": "1", "vag|ADJ": "1", "äntligen|ADV": "1", "vänster|ADJ": "1", "ner (el. ned)|ADV": "1", "väcka|VERB": "1", "leta|VERB": "1", "häst|NOUN": "1", "kategori|NOUN": "1", "brittisk|ADJ": "1", "följd|NOUN": "1", "ed|NOUN": "1", "fred|NOUN": "1", "traditionell|ADJ": "1", "användning|NOUN": "1", "riskera|VERB": "1", "tappa|VERB": "1", "inkomst|NOUN": "1", "nöjd|ADJ": "1", "kläder|NOUN": "1", "spara|VERB": "1", "styrelse|NOUN": "1", "intervju|NOUN": "1", "starkt|ADV": "1", "slutligen|ADV": "1", "bit|NOUN": "1", "muslimsk|ADJ": "1", "vetenskaplig|ADJ": "1", "överens|ADV": "1", "framtida|ADJ": "1", "bevis|NOUN": "1", "fast|ADJ": "1", "sexuell|ADJ": "1", "exakt|ADV": "1", "arbetsmarknad|NOUN": "1", "underbar|ADJ": "1", "post|NOUN": "1", "extra|ADJ": "1", "offer|NOUN": "1", "sektor|NOUN": "1", "vinst|NOUN": "1", "England|PROPN": "1", "inflytande|NOUN": "1", "budskap|NOUN": "1", "klicka|VERB": "1", "tips|NOUN": "1", "världskrig|NOUN": "1", "med tanke på|ADP": "1", "självklar|ADJ": "1", "båt|NOUN": "1", "borta|ADV": "1", "regional|ADJ": "1", "framåt|ADV": "1", "karaktär|NOUN": "1", "skiva|NOUN": "1", "omkring|ADV": "1", "ansikte|NOUN": "1", "i början|ADP": "1", "aktivitet|NOUN": "1", "ost|NOUN": "1", "fängelse|NOUN": "1", "motsvarande|ADJ": "1", "synas|VERB": "1", "mor (el. moder, vardagl. morsa) |NOUN": "1", "an|PART": "1", "samman|PART": "1", "ända|ADV": "1", "ledamot|NOUN": "1", "i enlighet med|ADP": "1", "civil|ADJ": "1", "uppenbar|ADJ": "1", "skull|NOUN": "1", "arbetslöshet|NOUN": "1", "fysisk|ADJ": "1", "generation|NOUN": "1", "återigen|ADV": "1", "djup|ADJ": "1", "initiativ|NOUN": "1", "fastställa|VERB": "1", "parlament|NOUN": "1", "säsong|NOUN": "1", "levande|ADJ": "1", "tacka|VERB": "1", "hota|VERB": "1", "tusentals|ADV": "1", "eventuell|ADJ": "1", "pojke|NOUN": "1", "version|NOUN": "1", "existera|VERB": "1", "trött|ADJ": "1", "himmel|NOUN": "1", "reaktion|NOUN": "1", "dyr|ADJ": "1", "normal|ADJ": "2", "rikta|VERB": "2", "kurs|NOUN": "2", "påstående|NOUN": "2", "märklig|ADJ": "2", "öst|NOUN": "2", "affär|NOUN": "2", "tidigt|ADV": "2", "upplevelse|NOUN": "2", "riktning|NOUN": "2", "vetenskap|NOUN": "2", "avsnitt|NOUN": "2", "handel|NOUN": "2", "sträckning|NOUN": "2", "locka|VERB": "2", "redovisa|VERB": "2", "uttalande|NOUN": "2", "respektive|CCONJ": "2", "para|VERB": "2", "störa|VERB": "2", "ihåg|PART": "2", "någonstans (vardagl. nånstans)|ADV": "2", "respekt|NOUN": "2", "rapportera|VERB": "2", "knappt|ADV": "2", "direkt|ADJ": "2", "enkelt|ADV": "2", "omständighet|NOUN": "2", "hänsyn|NOUN": "2", "ikväll (el. i kväll)|ADV": "2", "begära|VERB": "2", "rubrik|NOUN": "2", "producera|VERB": "2", "utsträckning|NOUN": "2", "anonym|ADJ": "2", "begå|VERB": "2", "bar|ADJ": "2", "institution|NOUN": "2", "förstöra|VERB": "2", "boll|NOUN": "2", "grunda|VERB": "2", "förbi|ADP": "2", "luft|NOUN": "2", "industri|NOUN": "2", "tåg|NOUN": "2", "skada|VERB": "2", "nordisk|ADJ": "2", "uppfylla|VERB": "2", "akta|VERB": "2", "förhandling|NOUN": "2", "syfta|VERB": "2", "bror (el. broder, vardagl. brorsa)|NOUN": "2", "byggnad|NOUN": "2", "hälft|NOUN": "2", "skrift|NOUN": "2", "ansvarig|ADJ": "2", "allmänhet|NOUN": "2", "orsaka|VERB": "2", "i slutet|ADP": "2", "israelisk|ADJ": "2", "drygt|ADV": "2", "lever|NOUN": "2", "bloggare|NOUN": "2", "tävling|NOUN": "2", "kommunikation|NOUN": "2", "kritisk|ADJ": "2", "plocka|VERB": "2", "patient|NOUN": "2", "sjunga|VERB": "2", "vakna|VERB": "2", "hälsa|NOUN": "2", "piratparti|NOUN": "2", "centrum|NOUN": "2", "otroligt|ADV": "2", "roligt|ADV": "2", "mörk|ADJ": "2", "träna|VERB": "2", "bord|NOUN": "2", "förrän|SCONJ": "2", "dansk|ADJ": "2", "vidta|VERB": "2", "reda|NOUN": "2", "mana|VERB": "2", "väljare|NOUN": "2", "uppmana|VERB": "2", "publik|NOUN": "2", "lida|VERB": "2", "motstånd|NOUN": "2", "lägenhet|NOUN": "2", "vänsterparti|NOUN": "2", "rädd|ADJ": "2", "användare|NOUN": "2", "inre|ADJ": "2", "avslöja|VERB": "2", "fiende|NOUN": "2", "lopp|NOUN": "2", "återvända|VERB": "2", "utmaning|NOUN": "2", "hopp|NOUN": "2", "konkurrens|NOUN": "2", "dröm|NOUN": "2", "detalj|NOUN": "2", "nedan|ADV": "2", "placera|VERB": "2", "litteratur|NOUN": "2", "ana|VERB": "2", "inställning|NOUN": "2", "armé|NOUN": "2", "lös|ADJ": "2", "pröva|VERB": "2", "egenskap|NOUN": "2", "rekommendera|VERB": "2", "liberal|ADJ": "2", "synpunkt|NOUN": "2", "undan|ADP": "2", "angående|ADP": "2", "unik|ADJ": "2", "präst|NOUN": "2", "webbplats|NOUN": "2", "bostad|NOUN": "2", "vardag|NOUN": "2", "gratis|ADV": "2", "återkomma|VERB": "2", "bevisa|VERB": "2", "anställd|NOUN": "2", "förbjuda|VERB": "2", "uttala|VERB": "2", "investering|NOUN": "2", "fira|VERB": "2", "försäljning|NOUN": "2", "populär|ADJ": "2", "klubb|NOUN": "2", "citat|NOUN": "2", "palestinier|NOUN": "2", "utrymme|NOUN": "2", "förr|ADV": "2", "svårt|ADV": "2", "stark|ADJ": "2", "påminna|VERB": "2", "aktör|NOUN": "2", "klassisk|ADJ": "2", "omkring|ADP": "2", "fokus|NOUN": "2", "officiell|ADJ": "2", "beröra|VERB": "2", "palestinsk|ADJ": "2", "ägare|NOUN": "2", "kapital|NOUN": "2", "relevant|ADJ": "2", "minister|NOUN": "2", "anpassa|VERB": "2", "glädje|NOUN": "2", "titel|NOUN": "2", "något|ADV": "2", "utgångspunkt|NOUN": "2", "nätverk|NOUN": "2", "scen|NOUN": "2", "nytta|NOUN": "2", "hållbar|ADJ": "2", "begränsa|VERB": "2", "sikte|NOUN": "2", "snygg|ADJ": "2", "kvinnlig|ADJ": "2", "som vanligt|ADV": "2", "avstånd|NOUN": "2", "fly|VERB": "2", "betydande|ADJ": "2", "skyldig|ADJ": "2", "i övrigt|ADV": "2", "inflation|NOUN": "2", "ben|NOUN": "2", "definition|NOUN": "2", "uppmärksamhet|NOUN": "2", "ladda|VERB": "2", "jul|NOUN": "2", "dåligt|ADV": "2", "kommunal|ADJ": "2", "passera|VERB": "2", "herre|NOUN": "2", "i fråga om|ADP": "2", "klimat|NOUN": "2", "var|PRON": "2", "topp|NOUN": "2", "troligen|ADV": "2", "kompis|NOUN": "2", "främja|VERB": "2", "landsting|NOUN": "2", "undersöka|VERB": "2", "kilometer (förk. km)|NOUN": "2", "reform|NOUN": "2", "testa|VERB": "2", "konkret|ADJ": "2", "rakt|ADV": "2", "uppenbarligen|ADV": "2", "desto|ADV": "2", "socialdemokratisk|ADJ": "2", "trupp|NOUN": "2", "vart|ADV": "2", "seger|NOUN": "2", "centerparti|NOUN": "2", "förlust|NOUN": "2", "själ|NOUN": "2", "öde|NOUN": "2", "mord|NOUN": "2", "dokument|NOUN": "2", "upphöra|VERB": "2", "folkparti|NOUN": "2", "kraftigt|ADV": "2", "middag|NOUN": "2", "reagera|VERB": "2", "hjärna|NOUN": "2", "kulturell|ADJ": "2", "södra|ADJ": "2", "fast|SCONJ": "2", "förtroende|NOUN": "2", "förordning|NOUN": "2", "upphovsrätt|NOUN": "2", "skuld|NOUN": "2", "professor|NOUN": "2", "inklusive|ADP": "2", "beskrivning|NOUN": "2", "lycka|NOUN": "2", "skrivning|NOUN": "2", "yrkande|NOUN": "2", "kär|ADJ": "2", "äng|NOUN": "2", "hänvisa|VERB": "2", "buss|NOUN": "2", "norra|ADJ": "2", "fullständigt|ADV": "2", "make|NOUN": "2", "antagligen|ADV": "2", "stil|NOUN": "2", "förbund|NOUN": "2", "tolkning|NOUN": "2", "utöver|ADP": "2", "syster (vardagl. syrra)|NOUN": "2", "berg|NOUN": "2", "motståndare|NOUN": "2", "höger|ADJ": "2", "praktisk|ADJ": "2", "beteende|NOUN": "2", "bud|NOUN": "2", "träning|NOUN": "2", "vare sig|CCONJ": "2", "äktenskap|NOUN": "2", "grov|ADJ": "2", "uppe|ADV": "2", "inslag|NOUN": "2", "förhindra|VERB": "2", "delning|NOUN": "2", "kapitalism|NOUN": "2", "bilaga|NOUN": "2", "tom|ADJ": "2", "invånare|NOUN": "2", "struktur|NOUN": "2", "politiskt|ADV": "2", "sjukhus|NOUN": "2", "mer eller mindre|ADV": "2", "främsta|ADJ": "2", "djupt|ADV": "2", "visning|NOUN": "2", "korrekt|ADJ": "2", "bäst|ADV": "2", "gentemot|ADP": "2", "tack vare|ADP": "2", "aspekt|NOUN": "2", "godkänna|VERB": "2", "felaktig|ADJ": "2", "dialog|NOUN": "2", "oro|NOUN": "2", "vägg|NOUN": "2", "kinesisk|ADJ": "2", "ständig|ADJ": "2", "tema|NOUN": "2", "helhet|NOUN": "2", "satsning|NOUN": "2", "statistik|NOUN": "2", "beräkna|VERB": "2", "resonemang|NOUN": "2", "förbud|NOUN": "2", "dollar|NOUN": "2", "längs|ADP": "2", "fixa|VERB": "2", "kollega|NOUN": "2", "inträffa|VERB": "2", "sjukvård|NOUN": "2", "överleva|VERB": "2", "sannolikt|ADV": "2", "i första hand|ADV": "2", "meddelande|NOUN": "2", "näringsliv|NOUN": "2", "låna|VERB": "2", "förståelse|NOUN": "2", "möjligen|ADV": "2", "fisk|NOUN": "2", "konsument|NOUN": "2", "framhålla|VERB": "2", "storlek|NOUN": "2", "telefon|NOUN": "2", "kön|NOUN": "2", "slut|PART": "2", "laga|VERB": "2", "roman|NOUN": "2", "lån|NOUN": "2", "likna|VERB": "2", "lita|VERB": "2", "säng|NOUN": "2", "rädsla|NOUN": "2", "övertygad|ADJ": "2", "skit|NOUN": "2", "tänkande|NOUN": "2", "arm|NOUN": "2", "bruk|NOUN": "2", "radio|NOUN": "2", "granska|VERB": "2", "i synnerhet|ADV": "2", "bekräfta|VERB": "2", "väder|NOUN": "2", "hinder|NOUN": "2", "förut|ADV": "2", "personligen|ADV": "2", "bana|NOUN": "2", "reklam|NOUN": "2", "trafik|NOUN": "2", "ärlig|ADJ": "2", "allting|PRON": "2", "artist|NOUN": "2", "bröd|NOUN": "2", "huruvida|SCONJ": "2", "utsatt|ADJ": "2", "butik|NOUN": "2", "ytterst|ADV": "2", "förbli|VERB": "2", "tråkig|ADJ": "2", "hemlig|ADJ": "2", "andlig|ADJ": "2", "beträffande|ADP": "2", "vänster|NOUN": "2", "fartyg|NOUN": "2", "flyga|VERB": "2", "gifta|VERB": "2", "snäll|ADJ": "2", "ränta|NOUN": "2", "proposition|NOUN": "2", "svårighet|NOUN": "2", "fart|NOUN": "2", "tant|NOUN": "2", "berörd|ADJ": "2", "avsikt|NOUN": "2", "frisk|ADJ": "2", "opposition|NOUN": "2", "härlig|ADJ": "2", "intryck|NOUN": "2", "visa|NOUN": "2", "duktig|ADJ": "2", "ideologi|NOUN": "2", "representant|NOUN": "2", "tack|NOUN": "2", "engagemang|NOUN": "2", "finsk|ADJ": "2", "bekant|ADJ": "2", "överallt|ADV": "2", "gäng|NOUN": "2", "träda|VERB": "2", "sjunka|VERB": "2", "föremål|NOUN": "2", "vad|ADV": "2", "attack|NOUN": "2", "falsk|ADJ": "2", "representera|VERB": "2", "miljöparti|NOUN": "2", "avgift|NOUN": "2", "normalt|ADV": "2", "motsvara|VERB": "2", "i allmänhet|ADV": "2", "översättning|NOUN": "2", "seriös|ADJ": "2", "omedelbart|ADV": "2", "kraftig|ADJ": "2", "uppskatta|VERB": "2", "kommitté|NOUN": "2", "blanda|VERB": "2", "blod|NOUN": "2", "högskola|NOUN": "2", "fritt|ADV": "2", "integritet|NOUN": "2", "hår|NOUN": "2", "organ|NOUN": "2", "lycklig|ADJ": "2", "misstag|NOUN": "2", "kvar|ADV": "2", "träd|NOUN": "2", "tak|NOUN": "2", "straff|NOUN": "2", "perfekt|ADJ": "2", "överenskommelse|NOUN": "2", "kampanj|NOUN": "2", "grej|NOUN": "2", "åstadkomma|VERB": "2", "budget|NOUN": "2", "rygg|NOUN": "2", "gott|ADV": "2", "press|NOUN": "2", "digital|ADJ": "2", "framstå|VERB": "2", "verktyg|NOUN": "2", "beroende på|ADP": "2", "betyg|NOUN": "2", "detsamma|PRON": "2", "start|NOUN": "2", "leverera|VERB": "2", "kompetens|NOUN": "2", "var och en|PRON": "2", "långsiktig|ADJ": "2", "vinter|NOUN": "2", "gripa|VERB": "2", "skyldighet|NOUN": "2", "evig|ADJ": "2", "företrädare|NOUN": "2", "etnisk|ADJ": "2", "med andra ord|ADV": "2", "njuta|VERB": "2", "posta|VERB": "2", "runda|VERB": "2", "för|CCONJ": "2", "bereda|VERB": "2", "uppmärksamma|VERB": "2", "arbetslös|ADJ": "2", "yta|NOUN": "2", "skratta|VERB": "2", "underlätta|VERB": "2", "föreligga|VERB": "2", "tillämpning|NOUN": "2", "garantera|VERB": "2", "jakt|NOUN": "2", "utse|VERB": "2", "blick|NOUN": "2", "svenska|NOUN": "2", "konferens|NOUN": "2", "framföra|VERB": "2", "runt|ADV": "2", "specifik|ADJ": "2", "varg|NOUN": "2", "kanal|NOUN": "2", "klok|ADJ": "2", "regim|NOUN": "2", "utöva|VERB": "2", "fokusera|VERB": "2", "belopp|NOUN": "2", "bransch|NOUN": "2", "sekund|NOUN": "2", "reda|VERB": "2", "torde|AUX": "2", "färdig|ADJ": "2", "ordna|VERB": "2", "närma|VERB": "2", "vind|NOUN": "2", "gård|NOUN": "2", "mitt|NOUN": "2", "framgångsrik|ADJ": "2", "identitet|NOUN": "2", "sång|NOUN": "2", "närma sig|VERB": "2", "skrika|VERB": "2", "tidpunkt|NOUN": "2", "avskaffa|VERB": "2", "samband|NOUN": "2", "lugn|ADJ": "2", "uppge|VERB": "2", "deltagare|NOUN": "2", "ursprung|NOUN": "2", "bestämd|ADJ": "2", "insikt|NOUN": "2", "forum|NOUN": "2", "kort|NOUN": "2", "statsminister|NOUN": "2", "annorlunda|ADJ": "2", "definiera|VERB": "2", "fönster|NOUN": "2", "get|NOUN": "2", "likhet|NOUN": "2", "ljud|NOUN": "2", "beställa|VERB": "2", "synd|NOUN": "2", "papper|NOUN": "2", "fara|NOUN": "2", "definitivt|ADV": "2", "omfattning|NOUN": "2", "bevara|VERB": "2", "väga|VERB": "2", "fenomen|NOUN": "2", "riktlinje|NOUN": "2", "profet|NOUN": "2", "decennium|NOUN": "2", "i stort sett|ADV": "2", "inriktning|NOUN": "2", "misslyckas|VERB": "2", "ram|NOUN": "2", "finansiera|VERB": "2", "hotell|NOUN": "2", "kristendom|NOUN": "2", "dess|ADV": "2", "i förhållande till|ADP": "2", "klaga|VERB": "2", "skatta|VERB": "2", "upprätta|VERB": "2", "förhoppningsvis|ADV": "2", "gynna|VERB": "2", "ifall|SCONJ": "2", "oberoende|ADJ": "2", "leka|VERB": "2", "märke|NOUN": "2", "snö|NOUN": "2", "upprepa|VERB": "2", "undervisning|NOUN": "2", "kött|NOUN": "2", "förutsätta|VERB": "2", "replik|NOUN": "2", "koppling|NOUN": "2", "snitt|NOUN": "2", "engelska|NOUN": "2", "överhuvudtaget|ADV": "2", "sysselsättning|NOUN": "2", "besked|NOUN": "2", "lätta|VERB": "2", "oavsett|ADV": "2", "avseende|NOUN": "2", "okänd|ADJ": "2", "katolsk|ADJ": "2", "ropa|VERB": "2", "bekämpa|VERB": "2", "synd|ADV": "2", "genast|ADV": "2", "sjö|NOUN": "2", "så småningom (el. småningom)|ADV": "2", "logisk|ADJ": "2", "inom ramen för|ADP": "2", "kaffe|NOUN": "2", "förstärka|VERB": "2", "euro|NOUN": "2", "mänsklighet|NOUN": "2", "nere|ADV": "2", "betona|VERB": "2", "expert|NOUN": "2", "fildelning|NOUN": "2", "olja|NOUN": "2", "förbereda|VERB": "2", "förfarande|NOUN": "2", "trygghet|NOUN": "2", "konstnär|NOUN": "2", "i själva verket|ADV": "2", "norsk|ADJ": "2", "i fråga (el. ifråga)|ADV": "2", "stjärna|NOUN": "2", "tyg|NOUN": "2", "läsning|NOUN": "2", "blå|ADJ": "2", "fotboll|NOUN": "2", "flykting|NOUN": "2", "koppla|VERB": "2", "forma|VERB": "2", "bibel|NOUN": "2", "förresten|ADV": "2", "samarbeta|VERB": "2", "slänga|VERB": "2", "ögonblick|NOUN": "2", "neka|VERB": "2", "extra|ADV": "2", "arbetsplats|NOUN": "2", "lokal|NOUN": "2", "summa|NOUN": "2", "tillräcklig|ADJ": "2", "äcklig|ADJ": "2", "tona|VERB": "2", "tendens|NOUN": "2", "på så sätt|ADV": "2", "restaurang|NOUN": "2", "återstå|VERB": "2", "vila|VERB": "2", "extremt|ADV": "2", "kamera|NOUN": "2", "självständig|ADJ": "2", "socialistisk|ADJ": "2", "framställa|VERB": "2", "ända (el. ände)|NOUN": "2", "mångfald|NOUN": "2", "strand|NOUN": "2", "pension|NOUN": "2", "hem|ADV": "2", "diskriminering|NOUN": "2", "misstänka|VERB": "2", "utsläpp|NOUN": "2", "logga|VERB": "2", "medicin|NOUN": "2", "sport|NOUN": "2", "rättvisa|NOUN": "2", "eld|NOUN": "2", "individuell|ADJ": "2", "därifrån|ADV": "2", "ifrån|ADV": "2", "yttre|ADJ": "2", "arabisk|ADJ": "2", "erhålla|VERB": "2", "moralisk|ADJ": "2", "revolutionär|ADJ": "2", "egendom|NOUN": "2", "köp|NOUN": "2", "välfärd|NOUN": "2", "sticka|VERB": "2", "mäta|VERB": "2", "helvete|NOUN": "2", "tuff|ADJ": "2", "jordbruk|NOUN": "2", "sällskap|NOUN": "2", "medverka|VERB": "2", "arbetstagare|NOUN": "2", "fånga|VERB": "2", "blogga|VERB": "2", "terrorism|NOUN": "2", "fest|NOUN": "2", "ordentligt|ADV": "2", "väst|NOUN": "2", "sajt|NOUN": "2", "prova|VERB": "2", "prägla|VERB": "2", "dum|ADJ": "2", "övning|NOUN": "2", "jobbig|ADJ": "2", "måla|VERB": "2", "vin|NOUN": "2", "identifiera|VERB": "2", "rasism|NOUN": "2", "ståndpunkt|NOUN": "2", "granne|NOUN": "2", "rang|NOUN": "2", "resultera|VERB": "2", "karriär|NOUN": "2", "trend|NOUN": "2", "kontor|NOUN": "2", "jaga|VERB": "2", "yttrandefrihet|NOUN": "2", "fortsättning|NOUN": "2", "diverse|ADJ": "2", "stöta|VERB": "2", "förneka|VERB": "2", "väsentlig|ADJ": "2", "manlig|ADJ": "2", "demonstration|NOUN": "2", "färd|NOUN": "2", "efterfrågan|NOUN": "2", "kandidat|NOUN": "2", "upprätthålla|VERB": "2", "fördrag|NOUN": "2", "instrument|NOUN": "2", "analysera|VERB": "2", "främmande|ADJ": "2", "uppmuntra|VERB": "2", "genomförande|NOUN": "2", "konservativ|ADJ": "2", "attityd|NOUN": "2", "föreställning|NOUN": "2", "än|SCONJ": "2", "lyda|VERB": "2", "juridisk|ADJ": "2", "variant|NOUN": "2", "höjd|NOUN": "2", "utrikesminister|NOUN": "2", "gäst|NOUN": "2", "hustru|NOUN": "2", "vandring|NOUN": "2", "kontakta|VERB": "2", "mil|NOUN": "2", "kort|ADV": "2", "eventuellt (förk. ev.)|ADV": "2", "lära|NOUN": "2", "medge|VERB": "2", "ologisk|ADJ": "2", "alkohol|NOUN": "2", "invandring|NOUN": "2", "arbetarklass|NOUN": "2", "lögn|NOUN": "2", "yttrande|NOUN": "2", "tillfällig|ADJ": "2", "varav|ADV": "2", "doktor (förk. dr)|NOUN": "2", "olaglig|ADJ": "2", "gränsa|VERB": "2", "vision|NOUN": "2", "framöver|ADV": "2", "över|ADV": "2", "omgivning|NOUN": "2", "bistånd|NOUN": "2", "ansluta|VERB": "2", "bas|NOUN": "2", "fil|NOUN": "2", "föredra|VERB": "2", "hemma|PART": "2", "sönder|PART": "2", "etablerad|ADJ": "2", "välkomna|VERB": "2", "tillverka|VERB": "2", "ambition|NOUN": "2", "aktie|NOUN": "2", "anklaga|VERB": "2", "dygn|NOUN": "2", "förtjäna|VERB": "2", "hur som helst (el. hursomhelst)|ADV": "2", "norm|NOUN": "2", "osäker|ADJ": "2", "räkning|NOUN": "2", "republik|NOUN": "2", "rykte|NOUN": "2", "jämförelse|NOUN": "2", "avstå|VERB": "2", "ära|NOUN": "2", "länsstyrelse|NOUN": "2", "smart|ADJ": "2", "bibliotek|NOUN": "2", "diktatur|NOUN": "2", "variera|VERB": "2", "dominera|VERB": "2", "utreda|VERB": "2", "boende|NOUN": "2", "museum|NOUN": "2", "förvandla|VERB": "2", "påbörja|VERB": "2", "ursäkt|NOUN": "2", "vete|NOUN": "2", "organisera|VERB": "2", "kommunistisk|ADJ": "2", "öra|NOUN": "2", "aktivt|ADV": "2", "granskning|NOUN": "2", "balans|NOUN": "2", "mage|NOUN": "2", "teckna|VERB": "2", "arg|ADJ": "2", "säkra|VERB": "2", "lunch|NOUN": "2", "kommunist|NOUN": "2", "militär|NOUN": "2", "gåva|NOUN": "2", "för närvarande|ADV": "2", "alternativ|ADJ": "2", "befintlig|ADJ": "2", "hälsa|VERB": "2", "socialism|NOUN": "2", "ursprunglig|ADJ": "2", "anställning|NOUN": "2", "ansökan|NOUN": "2", "protest|NOUN": "2", "test|NOUN": "3", "anda|NOUN": "2", "galen|ADJ": "2", "katastrof|NOUN": "2", "hata|VERB": "2", "gissa|VERB": "2", "mur|NOUN": "2", "tjänsteman|NOUN": "2", "led|NOUN": "4", "beakta|VERB": "2", "till följd av|ADP": "2", "reglera|VERB": "2", "kristdemokrat|NOUN": "2", "flod|NOUN": "2", "talare|NOUN": "2", "mörker|NOUN": "2", "begränsning|NOUN": "2", "värme|NOUN": "2", "agerande|NOUN": "2", "minoritet|NOUN": "2", "etablera|VERB": "2", "dam|NOUN": "2", "spansk|ADJ": "2", "motiv|NOUN": "2", "olikhet|NOUN": "2", "rättslig|ADJ": "2", "utställning|NOUN": "2", "utomlands|ADV": "2", "huvudstad|NOUN": "2", "likt|ADV": "2", "terrorist|NOUN": "2", "besökare|NOUN": "2", "hushåll|NOUN": "2", "respektera|VERB": "2", "fullständig|ADJ": "2", "mäktig|ADJ": "2", "växande|ADJ": "2", "stabil|ADJ": "2", "förvaltning|NOUN": "2", "hat|NOUN": "2", "mönster|NOUN": "2", "nyss|ADV": "2", "varumärke|NOUN": "2", "fastighet|NOUN": "2", "inta|VERB": "2", "orolig|ADJ": "2", "rulla|VERB": "2", "moral|NOUN": "2", "motivera|VERB": "2", "myt|NOUN": "2", "noga|ADV": "2", "snacka|VERB": "2", "till sist|ADV": "2", "förmedla|VERB": "2", "hamn|NOUN": "2", "tillhandahålla|VERB": "2", "informera|VERB": "2", "karta|NOUN": "2", "utforma|VERB": "2", "konvention|NOUN": "2", "allt mer (el. alltmer)|ADV": "2", "koll|NOUN": "2", "längd|NOUN": "2", "medicinsk|ADJ": "2", "läggning|NOUN": "2", "kilogram (el. kilo; förk. kg)|NOUN": "2", "finansiering|NOUN": "2", "löfte|NOUN": "2", "mörda|VERB": "2", "anställd|ADJ": "2", "amerikan|NOUN": "2", "rit|NOUN": "2", "status|NOUN": "2", "biologisk|ADJ": "2", "dikt|NOUN": "2", "sko|NOUN": "2", "sträcka|VERB": "2", "medarbetare|NOUN": "2", "lust|NOUN": "2", "kassa|NOUN": "2", "flygplats|NOUN": "2", "tingsrätt|NOUN": "2", "avdelning|NOUN": "2", "säkerställa|VERB": "2", "åklagare|NOUN": "2", "lysa|VERB": "2", "lidande|NOUN": "2", "syna|VERB": "2", "standard|NOUN": "2", "olycka|NOUN": "2", "term|NOUN": "2", "maskin|NOUN": "2", "transport|NOUN": "2", "etisk|ADJ": "2", "fattigdom|NOUN": "2", "servera|VERB": "2", "intern|ADJ": "2", "trolig|ADJ": "2", "golv|NOUN": "2", "förmiddag (förk. fm.)|NOUN": "2", "statsråd|NOUN": "2", "inrätta|VERB": "2", "närhet|NOUN": "2", "semester|NOUN": "2", "därigenom|ADV": "2", "ras|NOUN": "2", "tysk|NOUN": "2", "favorit|NOUN": "2", "framsteg|NOUN": "2", "tillvaro|NOUN": "2", "faktisk|ADJ": "2", "stolt|ADJ": "2", "strax|ADV": "2", "strida|VERB": "2", "angelägen|ADJ": "2", "skylla|VERB": "2", "ont|ADV": "2", "engagera|VERB": "2", "beräkning|NOUN": "2", "välkommen|ADJ": "2", "ideologisk|ADJ": "2", "finger|NOUN": "2", "hål|NOUN": "2", "prövning|NOUN": "2", "vettig|ADJ": "2", "komplicerad|ADJ": "2", "sund|ADJ": "2", "domare|NOUN": "2", "frukt|NOUN": "2", "signal|NOUN": "2", "guld|NOUN": "2", "homosexuell|ADJ": "2", "brottslighet|NOUN": "2", "rejäl|ADJ": "2", "rättegång|NOUN": "2", "mått|NOUN": "2", "kammare|NOUN": "2", "nazist|NOUN": "2", "förefalla|VERB": "2", "efteråt|ADV": "2", "försäkring|NOUN": "2", "konung|NOUN": "2", "såklart|ADV": "2", "ändamål|NOUN": "2", "avsedd|ADJ": "2", "generell|ADJ": "2", "kommunism|NOUN": "2", "dölja|VERB": "2", "arab|NOUN": "2", "sträva|VERB": "2", "stämning|NOUN": "2", "torg|NOUN": "2", "planerad|ADJ": "2", "utrustning|NOUN": "2", "vandra|VERB": "2", "registrera|VERB": "2", "argumentera|VERB": "2", "kök|NOUN": "2", "uppgå|VERB": "2", "visst|INTJ": "2", "bön|NOUN": "2", "anläggning|NOUN": "2", "filosofi|NOUN": "2", "gråta|VERB": "2", "underlag|NOUN": "2", "typisk|ADJ": "2", "förespråka|VERB": "2", "smärta|NOUN": "2", "uppror|NOUN": "2", "strategisk|ADJ": "2", "symbol|NOUN": "2", "radikal|ADJ": "2", "VD (verkställande direktör)|NOUN": "2", "frid|NOUN": "2", "arbetskraft|NOUN": "2", "bevilja|VERB": "2", "rot|NOUN": "2", "förmå|VERB": "2", "rak|ADJ": "2", "formulera|VERB": "2", "jämställdhet|NOUN": "2", "existens|NOUN": "2", "bonde|NOUN": "2", "bränna|VERB": "2", "italiensk|ADJ": "2", "utgift|NOUN": "2", "förbättring|NOUN": "2", "föreställa|VERB": "2", "operation|NOUN": "2", "landa|VERB": "2", "service|NOUN": "2", "låsa|VERB": "2", "varna|VERB": "2", "anställa|VERB": "2", "förtryck|NOUN": "2", "varelse|NOUN": "2", "tyst|ADJ": "2", "bredvid|ADP": "2", "syssla|VERB": "2", "drömma|VERB": "2", "evangelium|NOUN": "2", "planet|NOUN": "2", "organiserad|ADJ": "2", "fält|NOUN": "2", "omröstning|NOUN": "2", "psykisk|ADJ": "2", "fåtal|NOUN": "2", "öppet|ADV": "2", "överväga|VERB": "2", "stopp|NOUN": "2", "tråd|NOUN": "2", "prov|NOUN": "2", "sinne|NOUN": "2", "sorg|NOUN": "2", "ensamt|ADV": "2", "gemensamt|ADV": "2", "bort|ADV": "2", "kommersiell|ADJ": "2", "före detta (förk. f.d., f d)|ADV": "2", "sist|ADV": "2", "i huvudsak|ADV": "2", "lämpa sig|VERB": "2", "annorlunda|ADV": "2", "lura|VERB": "2", "förvisso|ADV": "2", "övervakning|NOUN": "2", "pågående|ADJ": "2", "utvärdering|NOUN": "2", "trygg|ADJ": "2", "arv|NOUN": "2", "seminarium|NOUN": "2", "besvara|VERB": "2", "övergrepp|NOUN": "2", "pass|NOUN": "2", "ljuga|VERB": "2", "uppdatering|NOUN": "2", "grekisk|ADJ": "2", "närvaro|NOUN": "2", "tidskrift|NOUN": "2", "infrastruktur|NOUN": "2", "biskop|NOUN": "2", "läger|NOUN": "2", "mer och mer|ADV": "2", "adress|NOUN": "2", "efterhand|ADV": "2", "förvånad|ADJ": "2", "ovanlig|ADJ": "2", "jävla (el. djävla)|ADJ": "2", "kontrakt|NOUN": "2", "skild|ADJ": "2", "daglig|ADJ": "2", "penningpolitik|NOUN": "2", "röstning|NOUN": "2", "lugnt|ADV": "2", "video|NOUN": "2", "med hänsyn till|ADP": "2", "översätta|VERB": "2", "fågel|NOUN": "2", "inkludera|VERB": "2", "era|NOUN": "2", "rörande|ADP": "2", "förena|VERB": "2", "ledig|ADJ": "2", "kärnkraft|NOUN": "2", "onödig|ADJ": "2", "ryss|NOUN": "2", "känslig|ADJ": "2", "smak|NOUN": "2", "order|NOUN": "2", "avancerad|ADJ": "2", "deltagande|NOUN": "2", "nämnd|NOUN": "2", "absolut|ADJ": "2", "israel|NOUN": "2", "prioritera|VERB": "2", "tillägga|VERB": "2", "blåsa|VERB": "2", "trädgård|NOUN": "2", "kors|NOUN": "2", "nyfiken|ADJ": "2", "kombination|NOUN": "2", "mod|NOUN": "2", "landskap|NOUN": "2", "överlämna|VERB": "2", "vinnare|NOUN": "2", "oskyldig|ADJ": "2", "fastna|VERB": "2", "förväntning|NOUN": "2", "temperatur|NOUN": "2", "övergripande|ADJ": "2", "motverka|VERB": "2", "våldsam|ADJ": "2", "fack|NOUN": "2", "komplettera|VERB": "2", "protokoll|NOUN": "2", "webb (el. web)|NOUN": "2", "bota|VERB": "2", "förlag|NOUN": "2", "bege sig|VERB": "2", "konsumtion|NOUN": "2", "värdefull|ADJ": "2", "kost|NOUN": "2", "godkänd|ADJ": "2", "datum|NOUN": "2", "därtill|ADV": "2", "recension|NOUN": "2", "till|ADV": "2", "omsorg|NOUN": "2", "kriterium|NOUN": "2", "fånge|NOUN": "2", "extrem|ADJ": "2", "förbindelse|NOUN": "2", "angrepp|NOUN": "2", "lansera|VERB": "2", "saga|NOUN": "2", "basera|VERB": "2", "cykel|NOUN": "2", "design|NOUN": "2", "frivillig|ADJ": "2", "med anledning av|ADP": "2", "västra|ADJ": "2", "påverkan|NOUN": "2", "verkan|NOUN": "2", "ful|ADJ": "2", "kongress|NOUN": "2", "skära|VERB": "2", "testamente|NOUN": "2", "gul|ADJ": "2", "skriftlig|ADJ": "2", "våg|NOUN": "2", "årlig|ADJ": "2", "reservation|NOUN": "2", "rättvis|ADJ": "2", "yrke|NOUN": "2", "århundrade|NOUN": "2", "anslag|NOUN": "2", "drog|NOUN": "2", "gömma|VERB": "2", "äkta|ADJ": "2", "intellektuell|ADJ": "2", "kejsare|NOUN": "2", "planering|NOUN": "2", "släkt|NOUN": "2", "drottning|NOUN": "2", "uppträda|VERB": "2", "övergå|VERB": "2", "het|ADJ": "2", "läkemedel|NOUN": "2", "utformning|NOUN": "2", "elektronisk|ADJ": "2", "obligatorisk|ADJ": "2", "investera|VERB": "2", "fond|NOUN": "2", "dubbel|ADJ": "2", "uppkomma|VERB": "2", "somna|VERB": "2", "ställningstagande|NOUN": "2", "utesluta|VERB": "2", "frukost|NOUN": "2", "förhoppning|NOUN": "2", "facklig|ADJ": "2", "prognos|NOUN": "2", "sannolikhet|NOUN": "2", "advokat|NOUN": "2", "kapitalistisk|ADJ": "2", "tveksam|ADJ": "2", "anlända|VERB": "2", "regn|NOUN": "2", "röja|VERB": "2", "motsats|NOUN": "2", "referens|NOUN": "2", "fabrik|NOUN": "2", "i och för sig|ADV": "2", "japansk|ADJ": "2", "plus|ADV": "2", "marknadsföring|NOUN": "2", "rena|VERB": "2", "innebörd|NOUN": "2", "stjäla|VERB": "2", "online|ADV": "2", "omgång|NOUN": "2", "protestera|VERB": "2", "tillkomma|VERB": "2", "bemöta|VERB": "2", "tränga|VERB": "2", "bestående|ADJ": "2", "blomma|NOUN": "2", "överföra|VERB": "2", "solidaritet|NOUN": "2", "lydelse|NOUN": "2", "annons|NOUN": "2", "riksdagsledamot|NOUN": "2", "brinna|VERB": "2", "rinna|VERB": "2", "gärning|NOUN": "2", "samverkan|NOUN": "2", "rymma|VERB": "2", "blogginlägg|NOUN": "2", "sammanfatta|VERB": "2", "östra|ADJ": "2", "dröja|VERB": "2", "avbryta|VERB": "2", "gräva|VERB": "2", "stryka|VERB": "2", "kreativ|ADJ": "2", "till dess|ADV": "2", "intensiv|ADJ": "2", "sålunda|ADV": "2", "roa|VERB": "2", "understryka|VERB": "2", "glas|NOUN": "2", "album|NOUN": "2", "territorium|NOUN": "2", "möjliggöra|VERB": "2", "fördelning|NOUN": "2", "folkomröstning|NOUN": "2", "skede|NOUN": "2", "markera|VERB": "2", "skaka|VERB": "2", "sten|NOUN": "2", "vagn|NOUN": "2", "värna|VERB": "2", "hemsk|ADJ": "2", "kriminell|ADJ": "2", "saklig|ADJ": "2", "närvarande|ADJ": "2", "automatiskt|ADV": "2", "skämma|VERB": "2", "vittna|VERB": "2", "spendera|VERB": "2", "ansvara|VERB": "2", "ledarskap|NOUN": "2", "trivas|VERB": "2", "figur|NOUN": "2", "bygd|NOUN": "2", "spridning|NOUN": "2", "lyckad|ADJ": "2", "le|VERB": "2", "betalning|NOUN": "2", "oroa|VERB": "2", "lov|NOUN": "2", "motsatt|ADJ": "2", "knyta|VERB": "2", "från och med|ADP": "2", "rekommendation|NOUN": "2", "ansträngning|NOUN": "2", "institut|NOUN": "2", "kritiker|NOUN": "2", "övre|ADJ": "2", "moderat|ADJ": "2", "data|NOUN": "2", "hörn|NOUN": "2", "inhemsk|ADJ": "2", "öl|NOUN": "2", "ängel|NOUN": "2", "blott|ADV": "2", "förhålla sig|VERB": "2", "förhålla|VERB": "2", "park|NOUN": "2", "regelverk|NOUN": "2", "nackdel|NOUN": "2", "vittne|NOUN": "2", "ljus|ADJ": "2", "medvetet|ADV": "2", "gas|NOUN": "2", "tipsa|VERB": "2", "våldtäkt|NOUN": "2", "boka|VERB": "2", "sådan här (vardagl. sån här)|DET": "2", "ekologisk|ADJ": "2", "återfinna|VERB": "2", "huvudsakligen|ADV": "2", "överge|VERB": "2", "ockupation|NOUN": "2", "likaså|ADV": "2", "bringa|VERB": "2", "hylla|VERB": "2", "sammanfattning|NOUN": "2", "liberal|NOUN": "2", "graf|NOUN": "2", "slott|NOUN": "2", "anspråk|NOUN": "2", "motsättning|NOUN": "2", "byte|NOUN": "2", "logik|NOUN": "2", "resonera|VERB": "2", "tempel|NOUN": "2", "krönika|NOUN": "2", "tillbringa|VERB": "2", "kopia|NOUN": "2", "instans|NOUN": "2", "företagare|NOUN": "2", "medlemskap|NOUN": "2", "egentlig|ADJ": "2", "landsbygd|NOUN": "2", "integration|NOUN": "2", "gest|NOUN": "2", "tyst|ADV": "2", "längta|VERB": "2", "föreskrift|NOUN": "2", "generellt|ADV": "2", "konto|NOUN": "2", "ju|CCONJ": "2", "tämligen|ADV": "2", "då och då|ADV": "2", "ryka|VERB": "2", "reglering|NOUN": "2", "misstänkt|ADJ": "2", "paket|NOUN": "2", "bete sig|VERB": "2", "kollektiv|ADJ": "2", "fotograf|NOUN": "2", "vänlig|ADJ": "2", "hemlighet|NOUN": "2", "administrativ|ADJ": "2", "dansa|VERB": "2", "tillägg|NOUN": "2", "fordon|NOUN": "2", "nöja sig|VERB": "2", "kliva|VERB": "2", "bro|NOUN": "2", "mandat|NOUN": "2", "inledning|NOUN": "2", "införande|NOUN": "2", "antyda|VERB": "2", "innefatta|VERB": "2", "kommunicera|VERB": "2", "praktiskt|ADV": "2", "förmån|NOUN": "2", "motivering|NOUN": "2", "tystnad|NOUN": "2", "valuta|NOUN": "2", "genomgå|VERB": "2", "nåd|NOUN": "2", "redaktion|NOUN": "2", "extern|ADJ": "2", "sfär|NOUN": "2", "flygplan|NOUN": "2", "kamrat|NOUN": "2", "premiärminister|NOUN": "2", "botten|NOUN": "2", "västerländsk|ADJ": "2", "skala|NOUN": "2", "utsikt|NOUN": "2", "besegra|VERB": "2", "utfärda|VERB": "2", "stimulera|VERB": "2", "kraftfull|ADJ": "2", "utöka|VERB": "2", "angripa|VERB": "2", "utseende|NOUN": "2", "promenad|NOUN": "2", "universum|NOUN": "2", "vanligtvis|ADV": "2", "pensionär|NOUN": "2", "redo|ADJ": "2", "järnväg|NOUN": "2", "jämn|ADJ": "2", "utbyte|NOUN": "2", "öppenhet|NOUN": "2", "grundval|NOUN": "2", "attackera|VERB": "2", "slita|VERB": "2", "förskola|NOUN": "2", "föregående|ADJ": "2", "föreskriva|VERB": "2", "inspiration|NOUN": "2", "anhängare|NOUN": "2", "hyra|VERB": "2", "kärna|NOUN": "2", "över huvud taget (el. överhuvudtaget)|ADV": "2", "löpa|VERB": "2", "blad|NOUN": "2", "gårdag|NOUN": "2", "tillföra|VERB": "2", "trovärdighet|NOUN": "2", "varv|NOUN": "2", "värdighet|NOUN": "2", "dans|NOUN": "2", "osäkerhet|NOUN": "2", "enstaka|ADJ": "2", "flyg|NOUN": "2", "vana|NOUN": "2", "spänning|NOUN": "2", "anfall|NOUN": "2", "utarbeta|VERB": "2", "skrämma|VERB": "2", "nyckel|NOUN": "2", "skribent|NOUN": "2", "garanti|NOUN": "2", "sakta|ADV": "2", "tillsätta|VERB": "2", "tvekan|NOUN": "2", "tand|NOUN": "2", "yrka|VERB": "2", "tacksam|ADJ": "2", "tävla|VERB": "2", "bortom|ADP": "2", "utbilda|VERB": "2", "hemland|NOUN": "2", "utav|ADP": "2", "avvisa|VERB": "2", "potentiell|ADJ": "2", "sovjetisk|ADJ": "2", "skepp|NOUN": "2", "utgång|NOUN": "2", "skrämmande|ADJ": "2", "omedelbar|ADJ": "2", "partner|NOUN": "2", "rejält|ADV": "2", "kapacitet|NOUN": "2", "genomsnitt|NOUN": "2", "värdig|ADJ": "2", "gymnasium|NOUN": "2", "umgås|VERB": "2", "knä|NOUN": "2", "element|NOUN": "2", "fredlig|ADJ": "2", "smal|ADJ": "2", "gubbe|NOUN": "2", "arrangera|VERB": "2", "skugga|NOUN": "2", "pressa|VERB": "2", "självständighet|NOUN": "2", "densamma|PRON": "2", "slutlig|ADJ": "2", "tvivel|NOUN": "2", "fälla|VERB": "2", "smaka|VERB": "2", "näst|ADV": "2", "utbud|NOUN": "2", "opinion|NOUN": "2", "värdera|VERB": "2", "allvarligt|ADV": "2", "formell|ADJ": "2", "dagligen|ADV": "2", "ursprungligen|ADV": "2", "vidare|ADJ": "2", "fördela|VERB": "2", "ovanligt|ADV": "2", "reducera|VERB": "2", "vanligt|ADV": "2", "skadestånd|NOUN": "2", "kopiera|VERB": "2", "övergång|NOUN": "2", "anhörig|ADJ": "2", "ångest|NOUN": "2", "vakt|NOUN": "2", "förhandla|VERB": "2", "koncentrera|VERB": "2", "tabell|NOUN": "2", "önskan|NOUN": "3", "konsert|NOUN": "3", "teckning|NOUN": "3", "avgå|VERB": "3", "grav|NOUN": "3", "agenda|NOUN": "3", "samfund|NOUN": "3", "krets|NOUN": "3", "kunglig|ADJ": "3", "anmälan|NOUN": "3", "inneha|VERB": "3", "soffa|NOUN": "3", "stabilitet|NOUN": "3", "förnuft|NOUN": "3", "därav|ADV": "3", "tredjedel|NOUN": "3", "ovanstående|ADJ": "3", "trovärdig|ADJ": "3", "strunta|VERB": "3", "akademisk|ADJ": "3", "permanent|ADJ": "3", "nyttig|ADJ": "3", "invändning|NOUN": "3", "våning|NOUN": "3", "långsamt|ADV": "3", "vild|ADJ": "3", "propaganda|NOUN": "3", "troende|ADJ": "3", "exemplar|NOUN": "3", "resolution|NOUN": "3", "ekonomiskt|ADV": "3", "därpå|ADV": "3", "formulering|NOUN": "3", "ihjäl|PART": "3", "såväl som|CCONJ": "3", "instämma|VERB": "3", "halvår|NOUN": "3", "debattera|VERB": "3", "idiot|NOUN": "3", "yttersta|ADJ": "3", "intill|ADP": "3", "torr|ADJ": "3", "söt|ADJ": "3", "socialist|NOUN": "3", "anordna|VERB": "3", "besviken|ADJ": "3", "lektion|NOUN": "3", "ledsen|ADJ": "3", "grattis|INTJ": "3", "sistnämnd|ADJ": "3", "tragisk|ADJ": "3", "teater|NOUN": "3", "försäkra|VERB": "3", "ideal|NOUN": "3", "vice|ADJ": "3", "hantering|NOUN": "3", "målsättning|NOUN": "3", "begripa|VERB": "3", "upphov|NOUN": "3", "kränka|VERB": "3", "i morse (el. imorse)|ADV": "3", "hals|NOUN": "3", "mån|NOUN": "3", "stam|NOUN": "3", "journalistik|NOUN": "3", "intäkt|NOUN": "3", "mjuk|ADJ": "3", "Bproper name (bruttonationalprodukt)|NOUN": "3", "grå|ADJ": "3", "profil|NOUN": "3", "krossa|VERB": "3", "partiledare|NOUN": "3", "centimeter (förk. cm)|NOUN": "3", "övertyga|VERB": "3", "romersk|ADJ": "3", "sörja|VERB": "3", "inspirera|VERB": "3", "övertygelse|NOUN": "3", "stackars|ADJ": "3", "sänkning|NOUN": "3", "potential|NOUN": "3", "antagande|NOUN": "3", "tilldela|VERB": "3", "biljett|NOUN": "3", "motsätta|VERB": "3", "komplex|ADJ": "3", "skadad|ADJ": "3", "begäran|NOUN": "3", "arena|NOUN": "3", "kust|NOUN": "3", "åtal|NOUN": "3", "dimension|NOUN": "3", "internationellt|ADV": "3", "nationellt|ADV": "3", "hållning|NOUN": "3", "gen|NOUN": "3", "lugn|NOUN": "3", "döpa|VERB": "3", "fantasi|NOUN": "3", "spets|NOUN": "3", "avsätta|VERB": "3", "fundering|NOUN": "3", "kombinera|VERB": "3", "observera|VERB": "3", "intressera|VERB": "3", "uppåt|ADV": "3", "fas|NOUN": "3", "dop|NOUN": "3", "professionell|ADJ": "3", "klippa|VERB": "3", "trist|ADJ": "3", "ombord|ADV": "3", "sparka|VERB": "3", "klimatförändring|NOUN": "3", "undervisa|VERB": "3", "dåvarande|ADJ": "3", "varning|NOUN": "3", "ton|NOUN": "3", "tänkbar|ADJ": "3", "villig|ADJ": "3", "station|NOUN": "3", "släkting|NOUN": "3", "övrigt|ADV": "3", "giltig|ADJ": "3", "gudomlig|ADJ": "3", "objektiv|ADJ": "3", "brand|NOUN": "3", "meningslös|ADJ": "3", "yttra|VERB": "3", "minskning|NOUN": "3", "axel|NOUN": "3", "försämra|VERB": "3", "motor|NOUN": "3", "i och med|ADV": "3", "konstruktion|NOUN": "3", "arkiv|NOUN": "3", "äventyr|NOUN": "3", "oj|INTJ": "3", "Sverige|PROPN": "3", "humor|NOUN": "3", "like|NOUN": "3", "paragraf|NOUN": "3", "odla|VERB": "3", "erbjudande|NOUN": "3", "vidga|VERB": "3", "volym|NOUN": "3", "motsätta sig|VERB": "3", "missbruk|NOUN": "3", "utvidga|VERB": "3", "snarast|ADV": "3", "uppmaning|NOUN": "3", "kram|NOUN": "3", "intervjua|VERB": "3", "livsmedel|NOUN": "3", "anklagelse|NOUN": "3", "cykla|VERB": "3", "samordning|NOUN": "3", "dessvärre|ADV": "3", "oklar|ADJ": "3", "företeelse|NOUN": "3", "offra|VERB": "3", "lager|NOUN": "3", "arbetsliv|NOUN": "3", "lysande|ADJ": "3", "bränsle|NOUN": "3", "finanskris|NOUN": "3", "nödvändigtvis|ADV": "3", "gott om|ADV": "3", "medeltid|NOUN": "3", "strävan|NOUN": "3", "hastighet|NOUN": "3", "kö|NOUN": "3", "medvetande|NOUN": "3", "producent|NOUN": "3", "så pass|ADV": "3", "vetande|NOUN": "3", "i mitten av|ADP": "3", "dylik|ADJ": "3", "installera|VERB": "3", "utge|VERB": "3", "förberedelse|NOUN": "3", "fördom|NOUN": "3", "synnerligen|ADV": "3", "i närheten av|ADP": "3", "åtagande|NOUN": "3", "tillkännage|VERB": "3", "kaos|NOUN": "3", "mästare|NOUN": "3", "utmana|VERB": "3", "drift|NOUN": "3", "hundratal|NOUN": "3", "måne|NOUN": "3", "bita|VERB": "3", "blandad|ADJ": "3", "hjälte|NOUN": "3", "skänka|VERB": "3", "tillämplig|ADJ": "3", "betydelsefull|ADJ": "3", "synsätt|NOUN": "3", "ström|NOUN": "3", "förse|VERB": "3", "mätning|NOUN": "3", "massiv|ADJ": "3", "atmosfär|NOUN": "3", "mall|NOUN": "3", "personlighet|NOUN": "3", "gren|NOUN": "3", "väldig|ADJ": "3", "effektivt|ADV": "3", "vanligen|ADV": "3", "koncept|NOUN": "3", "välkänd|ADJ": "3", "förebild|NOUN": "3", "uppenbart|ADV": "3", "recept|NOUN": "3", "föreläsning|NOUN": "3", "antisemitism|NOUN": "3", "geografisk|ADJ": "3", "grafisk|ADJ": "3", "upplysning|NOUN": "3", "general|NOUN": "3", "administration|NOUN": "3", "bröst|NOUN": "3", "tills|ADP": "3", "patent|NOUN": "3", "befogenhet|NOUN": "3", "skarp|ADJ": "3", "islamisk|ADJ": "3", "vem som helst|PRON": "3", "förverkliga|VERB": "3", "prioritering|NOUN": "3", "vistas|VERB": "3", "regelbundet|ADV": "3", "depression|NOUN": "3", "effektivitet|NOUN": "3", "inne|PART": "3", "likväl|ADV": "3", "blandning|NOUN": "3", "datera|VERB": "3", "final|NOUN": "3", "tjock|ADJ": "3", "erövra|VERB": "3", "höger|NOUN": "3", "sträcka|NOUN": "3", "vaka|VERB": "3", "polsk|ADJ": "3", "bomb|NOUN": "3", "tår|NOUN": "3", "fackförening|NOUN": "3", "utvald|ADJ": "3", "placering|NOUN": "3", "huvudsaklig|ADJ": "3", "avfall|NOUN": "3", "gigantisk|ADJ": "3", "väntan|NOUN": "3", "turnering|NOUN": "3", "uppvärmning|NOUN": "3", "djup|NOUN": "3", "praxis|NOUN": "3", "okej|INTJ": "3", "maximal (förk. max.)|ADJ": "3", "konstitution|NOUN": "3", "otrolig|ADJ": "3", "fruktansvärd|ADJ": "3", "straffa|VERB": "3", "sådär|ADV": "3", "nödvändighet|NOUN": "3", "medlemsland|NOUN": "3", "översyn|NOUN": "3", "blind|ADJ": "3", "front|NOUN": "3", "fördöma|VERB": "3", "synlig|ADJ": "3", "fint|ADV": "3", "skapelse|NOUN": "3", "rasa|VERB": "3", "verksam|ADJ": "3", "avlida|VERB": "3", "fullkomligt|ADV": "3", "teoretisk|ADJ": "3", "flyta|VERB": "3", "urval|NOUN": "3", "binda|VERB": "3", "fett|NOUN": "3", "erkännande|NOUN": "3", "hälsning|NOUN": "3", "idrott|NOUN": "3", "debattartikel|NOUN": "3", "belysa|VERB": "3", "emellan|ADP": "3", "övervaka|VERB": "3", "lagom|ADV": "3", "sömn|NOUN": "3", "proletariat|NOUN": "3", "önskemål|NOUN": "3", "förlåta|VERB": "3", "sammanlagt|ADV": "3", "slav|NOUN": "3", "näsa|NOUN": "3", "däribland|ADV": "3", "export|NOUN": "3", "nedgång|NOUN": "3", "vinkel|NOUN": "3", "experiment|NOUN": "3", "allierad|ADJ": "3", "arbetstid|NOUN": "3", "flagga|NOUN": "3", "uppdatera|VERB": "3", "block|NOUN": "3", "feminism|NOUN": "3", "skattebetalare|NOUN": "3", "globalisering|NOUN": "3", "miljontals|ADV": "3", "obehaglig|ADJ": "3", "ondska|NOUN": "3", "önskvärd|ADJ": "3", "anpassad|ADJ": "3", "mysig|ADJ": "3", "norr|NOUN": "3", "andning|NOUN": "3", "motta|VERB": "3", "utspela sig|VERB": "3", "exakt|ADJ": "3", "elit|NOUN": "3", "inverkan|NOUN": "3", "akut|ADJ": "3", "kvarstå|VERB": "3", "troligtvis|ADV": "3", "konkurs|NOUN": "3", "center|NOUN": "3", "än så länge|ADV": "3", "dramatisk|ADJ": "3", "låtsas|VERB": "3", "underlig|ADJ": "3", "förlängning|NOUN": "3", "segla|VERB": "3", "försiktig|ADJ": "3", "himla|ADV": "3", "inbördeskrig|NOUN": "3", "vid sidan av|ADP": "3", "grym|ADJ": "3", "tunn|ADJ": "3", "grundlag|NOUN": "3", "realistisk|ADJ": "3", "tvätta|VERB": "3", "enormt|ADV": "3", "litterär|ADJ": "3", "mobiltelefon|NOUN": "3", "dominerande|ADJ": "3", "framkomma|VERB": "3", "misshandel|NOUN": "3", "skildra|VERB": "3", "förbannad|ADJ": "3", "anpassning|NOUN": "3", "redaktör|NOUN": "3", "behörig|ADJ": "3", "last|NOUN": "3", "arbetarrörelse|NOUN": "3", "liberalism|NOUN": "3", "presentation|NOUN": "3", "stress|NOUN": "3", "försörja|VERB": "3", "objekt|NOUN": "3", "omslag|NOUN": "3", "absurd|ADJ": "3", "kvalificerad|ADJ": "3", "trappa|NOUN": "3", "offentligt|ADV": "3", "röka|VERB": "3", "valrörelse|NOUN": "3", "anfalla|VERB": "3", "rådande|ADJ": "3", "spåra|VERB": "3", "upplaga|NOUN": "3", "ordentlig|ADJ": "3", "klä (el. kläda)|VERB": "3", "ambassad|NOUN": "3", "konkurrera|VERB": "3", "ovanför|ADP": "3", "skämt|NOUN": "3", "tända|VERB": "3", "anslutning|NOUN": "3", "backa|VERB": "3", "loss|PART": "3", "samvete|NOUN": "3", "fastän|SCONJ": "3", "årtionde|NOUN": "3", "tomt|NOUN": "3", "avsevärt|ADV": "3", "rita|VERB": "3", "värt|ADV": "3", "register|NOUN": "3", "rörlighet|NOUN": "3", "ignorera|VERB": "3", "dold|ADJ": "3", "befria|VERB": "3", "först och främst|ADV": "3", "retorik|NOUN": "3", "leende|NOUN": "3", "olycklig|ADJ": "3", "säkerligen|ADV": "3", "abort|NOUN": "3", "taktik|NOUN": "3", "beteckna|VERB": "3", "lärjunge|NOUN": "3", "stadga|NOUN": "3", "långsam|ADJ": "3", "oberoende av|ADP": "3", "utlänning|NOUN": "3", "spelning|NOUN": "3", "godkännande|NOUN": "3", "fet|ADJ": "3", "hovrätt|NOUN": "3", "tiotal|NOUN": "3", "skivbolag|NOUN": "3", "stycke|NOUN": "3", "tempo|NOUN": "3", "påve|NOUN": "3", "kant|NOUN": "3", "turist|NOUN": "3", "predika|VERB": "3", "reflektera|VERB": "3", "folkgrupp|NOUN": "3", "rektor|NOUN": "3", "klargöra|VERB": "3", "neutral|ADJ": "3", "laglig|ADJ": "3", "tendera|VERB": "3", "utrikespolitik|NOUN": "3", "glädja|VERB": "3", "rödgrön|ADJ": "3", "segra|VERB": "3", "inrikta|VERB": "3", "monopol|NOUN": "3", "konkurrent|NOUN": "3", "plattform|NOUN": "3", "skådespelare|NOUN": "3", "störning|NOUN": "3", "remissinstans|NOUN": "3", "rutin|NOUN": "3", "dal|NOUN": "3", "studio|NOUN": "3", "användbar|ADJ": "3", "lagförslag|NOUN": "3", "självfallet|ADV": "3", "ömsesidig|ADJ": "3", "förvåna|VERB": "3", "flaska|NOUN": "3", "packa|VERB": "3", "reportage|NOUN": "3", "skylt|NOUN": "3", "platta|NOUN": "3", "välsignelse|NOUN": "3", "cell|NOUN": "3", "i förväg|ADV": "3", "kopp|NOUN": "3", "bortse|VERB": "3", "etik|NOUN": "3", "mördare|NOUN": "3", "med stöd av|ADP": "3", "vid|ADJ": "3", "förintelse|NOUN": "3", "redogöra|VERB": "3", "auktoritet|NOUN": "3", "avslå|VERB": "3", "hud|NOUN": "3", "välstånd|NOUN": "3", "rättfärdig|ADJ": "3", "därvid|ADV": "3", "tillgodose|VERB": "3", "mental|ADJ": "3", "försvarsmakt|NOUN": "3", "kollektivavtal|NOUN": "3", "svaghet|NOUN": "3", "frågeställning|NOUN": "3", "motsvarighet|NOUN": "3", "slutändan|NOUN": "3", "bitter|ADJ": "3", "utanförskap|NOUN": "3", "åtskillig|ADJ": "3", "koldioxid|NOUN": "3", "mässa|NOUN": "3", "rå|ADJ": "3", "tvivla|VERB": "3", "höjning|NOUN": "3", "forn|ADJ": "3", "konjunktur|NOUN": "3", "nöje|NOUN": "3", "attraktiv|ADJ": "3", "reflektion|NOUN": "3", "samråd|NOUN": "3", "afrikansk|ADJ": "3", "kontroversiell|ADJ": "3", "ruta|NOUN": "3", "folklig|ADJ": "3", "framträda|VERB": "3", "vis|ADJ": "3", "förlänga|VERB": "3", "spegla|VERB": "3", "frånvaro|NOUN": "3", "symptom (el. symtom)|NOUN": "3", "bokstav|NOUN": "3", "webbläsare|NOUN": "3", "skrivelse|NOUN": "3", "barndom|NOUN": "3", "usel|ADJ": "3", "folkmord|NOUN": "3", "till känna|ADV": "3", "arbetsuppgift|NOUN": "3", "illegal|ADJ": "3", "städa|VERB": "3", "uppvisa|VERB": "3", "väska|NOUN": "3", "ärligt|ADV": "3", "historiskt|ADV": "3", "upphovsman|NOUN": "3", "lock|NOUN": "3", "tes|NOUN": "3", "bekostnad|NOUN": "3", "info|NOUN": "3", "skadlig|ADJ": "3", "ansöka|VERB": "3", "industriell|ADJ": "3", "köpare|NOUN": "3", "börs|NOUN": "3", "beklaga|VERB": "3", "korruption|NOUN": "3", "uppföra|VERB": "3", "arbetsförmedling|NOUN": "3", "fria|VERB": "3", "britt|NOUN": "3", "kontinent|NOUN": "3", "låda|NOUN": "3", "bevaka|VERB": "3", "besparing|NOUN": "3", "redovisning|NOUN": "3", "variation|NOUN": "3", "detaljerad|ADJ": "3", "skratt|NOUN": "3", "naken|ADJ": "3", "byggande|NOUN": "3", "konstruktiv|ADJ": "3", "integrera|VERB": "3", "återkommande|ADJ": "3", "slump|NOUN": "3", "mottagare|NOUN": "3", "återgå|VERB": "3", "i likhet med|ADV": "3", "leverantör|NOUN": "3", "noll|NUM": "3", "storm|NOUN": "3", "pirat|NOUN": "3", "svänga|VERB": "3", "bifall|NOUN": "3", "instruktion|NOUN": "3", "upptagen|ADJ": "3", "paus|NOUN": "3", "rationell|ADJ": "3", "överstiga|VERB": "3", "delad|ADJ": "3", "skärpa|VERB": "3", "tillverkare|NOUN": "3", "imponerande|ADJ": "3", "följaktligen|ADV": "3", "innan|ADP": "3", "misstanke|NOUN": "3", "omdöme|NOUN": "3", "kod|NOUN": "3", "server|NOUN": "3", "magisk|ADJ": "3", "sträng|ADJ": "3", "vad som helst|ADV": "3", "dagbok|NOUN": "3", "radera|VERB": "3", "anknytning|NOUN": "3", "häromdagen|ADV": "3", "innovation|NOUN": "3", "gran|NOUN": "3", "uppföljning|NOUN": "3", "grabb|NOUN": "3", "frukta|VERB": "3", "tvist|NOUN": "3", "innan|ADV": "3", "van|ADJ": "3", "dubbelt|ADV": "3", "mild|ADJ": "3", "drivkraft|NOUN": "3", "tjänare|NOUN": "3", "nationalism|NOUN": "3", "moln|NOUN": "3", "ordförandeskap|NOUN": "3", "såvitt|SCONJ": "3", "mekanism|NOUN": "3", "minsann|ADV": "3", "vaccin|NOUN": "3", "filosof|NOUN": "3", "division|NOUN": "3", "belägen|ADJ": "3", "tåla|VERB": "3", "avdrag|NOUN": "3", "koloni|NOUN": "3", "sannerligen|ADV": "3", "till förmån för|ADP": "3", "cancer|NOUN": "3", "förföljelse|NOUN": "3", "byråkrati|NOUN": "3", "mobil|ADJ": "3", "tillsyn|NOUN": "3", "ett|PRON": "3", "sur|ADJ": "3", "nazism|NOUN": "3", "rösträtt|NOUN": "3", "somlig|PRON": "3", "utredare|NOUN": "3", "stadium|NOUN": "3", "dagis|NOUN": "3", "färsk|ADJ": "3", "positivt|ADV": "3", "livsstil|NOUN": "3", "pressmeddelande|NOUN": "3", "klyfta|NOUN": "3", "skapande|NOUN": "3", "inlagd|ADJ": "3", "konstnärlig|ADJ": "3", "pinsam|ADJ": "3", "löpande|ADJ": "3", "konstant|ADJ": "3", "åberopa|VERB": "3", "arrangemang|NOUN": "3", "avslutad|ADJ": "3", "varifrån|ADV": "3", "jurist|NOUN": "3", "lagra|VERB": "3", "påtaglig|ADJ": "3", "tillgänglighet|NOUN": "3", "pedagogisk|ADJ": "3", "skita|VERB": "3", "kärnvapen|NOUN": "3", "plikt|NOUN": "3", "företräda|VERB": "3", "mjölk|NOUN": "3", "policy|NOUN": "3", "ångra|VERB": "3", "apostel|NOUN": "3", "ingripa|VERB": "3", "tröttna|VERB": "3", "utvidgning|NOUN": "3", "kvarter|NOUN": "3", "flexibel|ADJ": "3", "motionär|NOUN": "3", "ideell|ADJ": "3", "insyn|NOUN": "3", "bosatt|ADJ": "3", "filosofisk|ADJ": "3", "inspelning|NOUN": "3", "reell|ADJ": "3", "generera|VERB": "3", "krypa|VERB": "3", "kränkning|NOUN": "3", "trogen|ADJ": "3", "underteckna|VERB": "3", "stilla|ADV": "3", "invasion|NOUN": "3", "enhetlig|ADJ": "3", "not|NOUN": "3", "förebygga|VERB": "3", "lukta|VERB": "3", "humanitär|ADJ": "3", "intelligent|ADJ": "3", "besvär|NOUN": "3", "flotta|NOUN": "3", "turkisk|ADJ": "3", "mandatperiod|NOUN": "3", "civilisation|NOUN": "3", "ursäkta|VERB": "3", "demonstrera|VERB": "3", "godta|VERB": "3", "andas|VERB": "3", "böter|NOUN": "3", "lärdom|NOUN": "3", "kyla|NOUN": "3", "ordinarie|ADJ": "3", "delegation|NOUN": "3", "suga|VERB": "3", "tränare|NOUN": "3", "användande|NOUN": "3", "arbetsgrupp|NOUN": "3", "operatör|NOUN": "3", "reporter|NOUN": "3", "tortyr|NOUN": "3", "kapten|NOUN": "3", "forska|VERB": "3", "avkastning|NOUN": "3", "genomsnittlig|ADJ": "3", "jägare|NOUN": "3", "makthavare|NOUN": "3", "löjlig|ADJ": "3", "skönhet|NOUN": "3", "orimlig|ADJ": "3", "matematik|NOUN": "3", "officiellt|ADV": "3", "rensa|VERB": "3", "utvärdera|VERB": "3", "onekligen|ADV": "3", "tonåring|NOUN": "3", "dagsläge|NOUN": "3", "entreprenör|NOUN": "3", "kines|NOUN": "3", "blivande|ADJ": "3", "elände|NOUN": "3", "glida|VERB": "3", "stiftelse|NOUN": "3", "frivilligt|ADV": "3", "introducera|VERB": "3", "korrekt|ADV": "3", "villigt|ADV": "3", "friskola|NOUN": "3", "smula|NOUN": "3", "försvåra|VERB": "3", "kyrklig|ADJ": "3", "oväntad|ADJ": "3", "rikedom|NOUN": "3", "delstat|NOUN": "3", "gång på gång|ADV": "3", "illustrera|VERB": "3", "centralbank|NOUN": "3", "grannland|NOUN": "3", "rasist|NOUN": "3", "ägande|NOUN": "3", "förvirrad|ADJ": "3", "kredit|NOUN": "3", "rom|NOUN": "3", "storstad|NOUN": "3", "tveka|VERB": "3", "överföring|NOUN": "3", "katolik|NOUN": "3", "tät|ADJ": "3", "fotografi|NOUN": "3", "förare|NOUN": "3", "historiker|NOUN": "3", "misslyckande|NOUN": "3", "present|NOUN": "3", "dödsstraff|NOUN": "3", "evighet|NOUN": "3", "enighet|NOUN": "3", "torn|NOUN": "3", "stigande|ADJ": "3", "förkasta|VERB": "3", "humör|NOUN": "3", "hemskt|ADV": "3", "moment|NOUN": "3", "allihop (vardagl. allihopa)|PRON": "3", "fritid|NOUN": "3", "rapportering|NOUN": "3", "stöld|NOUN": "3", "konkurrenskraft|NOUN": "3", "psykologisk|ADJ": "3", "alternativt|ADV": "3", "direktör|NOUN": "3", "skeptisk|ADJ": "3", "bakåt|ADV": "3", "lapp|NOUN": "3", "anlita|VERB": "3", "avfärda|VERB": "3", "likadant|ADV": "3", "separat|ADJ": "3", "överensstämma|VERB": "3", "finansminister|NOUN": "3", "format|NOUN": "3", "ogilla|VERB": "3", "omvandla|VERB": "3", "argumentation|NOUN": "3", "likadan|ADJ": "3", "tavla|NOUN": "3", "kännedom|NOUN": "3", "programvara|NOUN": "3", "skattesänkning|NOUN": "3", "jämlikhet|NOUN": "3", "chefredaktör|NOUN": "3", "säljare|NOUN": "3", "duga|VERB": "3", "negativt|ADV": "3", "arkitekt|NOUN": "3", "livad|ADJ": "3", "passagerare|NOUN": "3", "finans|NOUN": "3", "ekonom|NOUN": "3", "läsvärd|ADJ": "3", "obegriplig|ADJ": "3", "skam|NOUN": "3", "skicklig|ADJ": "3", "störta|VERB": "3", "överta|VERB": "3", "feminist|NOUN": "3", "orättvisa|NOUN": "3", "stadsdel|NOUN": "3", "årligen|ADV": "3", "utbyggnad|NOUN": "3", "beskattning|NOUN": "3", "återge|VERB": "3", "koka|VERB": "3", "taliban|NOUN": "3", "skara|NOUN": "3", "bröllop|NOUN": "3", "mormor|NOUN": "3", "pasta|NOUN": "3", "itu|PART": "3", "fan|NOUN": "3", "syskon|NOUN": "3", "tillverkning|NOUN": "3", "bunden|ADJ": "3", "gitarr|NOUN": "3", "diagnos|NOUN": "3", "häftig|ADJ": "3", "överklaga|VERB": "3", "strejk|NOUN": "3", "tvång|NOUN": "3", "dödsfall|NOUN": "3", "import|NOUN": "3", "formellt|ADV": "3", "rund|ADJ": "3", "sambo|NOUN": "3", "teknologi|NOUN": "3", "iransk|ADJ": "3", "någorlunda|ADV": "3", "genomgång|NOUN": "3", "grundskola|NOUN": "3", "framställning|NOUN": "3", "rådgivare|NOUN": "3", "vrida|VERB": "3", "behaglig|ADJ": "3", "fästa|VERB": "3", "målning|NOUN": "3", "underskott|NOUN": "3", "framme|ADV": "3", "imperium|NOUN": "3", "lönsam|ADJ": "3", "söder|NOUN": "3", "successivt|ADV": "3", "hänvisning|NOUN": "3", "konsekvent|ADV": "3", "isolerad|ADJ": "3", "handlingsplan|NOUN": "3", "tvåa|NOUN": "3", "häva|VERB": "3", "upphäva|VERB": "3", "färdighet|NOUN": "3", "självmord|NOUN": "3", "svärd|NOUN": "3", "stall|NOUN": "3", "styre|NOUN": "3", "fristående|ADJ": "3", "ilska|NOUN": "3", "dumt|ADJ": "3", "offentliggöra|VERB": "3", "privatperson|NOUN": "3", "kompensera|VERB": "3", "överraskning|NOUN": "3", "stängd|ADJ": "3", "tröja|NOUN": "3", "komponent|NOUN": "3", "festival|NOUN": "3", "lågkonjunktur|NOUN": "3", "återställa|VERB": "3", "skandal|NOUN": "3", "med hänvisning till|ADP": "3", "förutse|VERB": "3", "minst sagt|ADV": "3", "stötta|VERB": "3", "fantastiskt|ADV": "3", "karl|NOUN": "3", "aggressiv|ADJ": "3", "härmed|ADV": "3", "avsaknad|NOUN": "3", "kemisk|ADJ": "3", "saknad|NOUN": "3", "raket|NOUN": "3", "tunnelbana|NOUN": "3", "värma|VERB": "3", "kommunistparti|NOUN": "3", "marginal|NOUN": "3", "respektive|ADV": "3", "gravid|ADJ": "3", "kniv|NOUN": "3", "ramla|VERB": "3", "villa|NOUN": "3", "dryg|ADJ": "3", "lampa|NOUN": "3", "överdriven|ADJ": "3", "back|NOUN": "3", "kusin|NOUN": "3", "knapp|NOUN": "3", "skynda|VERB": "3", "privatliv|NOUN": "3", "toalett|NOUN": "3", "bada|VERB": "3", "lustig|ADJ": "3", "provins|NOUN": "3", "orättvis|ADJ": "3", "sexualitet|NOUN": "3", "upptäckt|NOUN": "3", "kreativitet|NOUN": "3", "lagråd|NOUN": "3", "malm|NOUN": "3", "referera|VERB": "3", "teologi|NOUN": "3", "arkitektur|NOUN": "3", "förvalta|VERB": "3", "rättsväsende|NOUN": "3", "lord|NOUN": "3", "poet|NOUN": "3", "stuga|NOUN": "3", "regna|VERB": "3", "spekulera|VERB": "3", "bonus|NOUN": "3", "längtan|NOUN": "3", "rymd|NOUN": "3", "fruktansvärt|ADV": "3", "bad|NOUN": "3", "förhör|NOUN": "3", "likvärdig|ADJ": "3", "upplösa|VERB": "3", "blockera|VERB": "3", "fröken|NOUN": "3", "hysa|VERB": "3", "klipp|NOUN": "3", "äganderätt|NOUN": "3", "akademi|NOUN": "3", "benämna|VERB": "3", "indisk|ADJ": "3", "rosa|ADJ": "3", "tycke|NOUN": "3", "avlägsen|ADJ": "3", "konstigt|ADV": "3", "marknadsekonomi|NOUN": "3", "uppta|VERB": "3", "utland|NOUN": "3", "erinra|VERB": "3", "finanser|NOUN": "3", "lärande|NOUN": "3", "råvara|NOUN": "3", "förenlig|ADJ": "3", "klättra|VERB": "3", "berättigad|ADJ": "3", "brottsling|NOUN": "3", "tillhörande|ADJ": "3", "delaktig|ADJ": "3", "rusa|VERB": "3", "änka|NOUN": "3", "plugga|VERB": "3", "prins|NOUN": "3", "mystisk|ADJ": "3", "same|NOUN": "3", "bar|NOUN": "3", "indirekt|ADV": "3", "webbsida|NOUN": "3", "avveckla|VERB": "3", "bygge|NOUN": "3", "föredrag|NOUN": "3", "bibehålla|VERB": "3", "näring|NOUN": "3", "poesi|NOUN": "3", "smyga|VERB": "3", "förort|NOUN": "3", "genetisk|ADJ": "3", "sorglig|ADJ": "3", "fransman|NOUN": "3", "genre|NOUN": "3", "lat|ADJ": "3", "lastbil|NOUN": "3", "vårda|VERB": "3", "lista|VERB": "3", "inledande|ADJ": "3", "debattör|NOUN": "3", "premiär|NOUN": "3", "redskap|NOUN": "3", "vila|NOUN": "3", "novell|NOUN": "3", "väsentligt|ADV": "3", "matte|NOUN": "3", "anförande|NOUN": "3", "hyra|NOUN": "3", "mogen|ADJ": "3", "osynlig|ADJ": "3", "besvärlig|ADJ": "3", "dansk|NOUN": "3", "överskott|NOUN": "3", "kompromiss|NOUN": "3", "uppskattning|NOUN": "3", "kvart|NOUN": "3", "spekulation|NOUN": "3", "urban|ADJ": "3", "begriplig|ADJ": "3", "träff|NOUN": "3", "flykt|NOUN": "3", "poker|NOUN": "3", "uppgörelse|NOUN": "3", "besvikelse|NOUN": "3", "gradvis|ADV": "3", "acceptabel|ADJ": "3", "lugna|VERB": "3", "skräck|NOUN": "3", "komplett|ADJ": "3", "norr om|ADP": "3", "förhållandevis|ADV": "3", "hugga|VERB": "3", "massmedium|NOUN": "3", "varpå|ADV": "3", "åtala|VERB": "3", "gris|NOUN": "3", "medverkan|NOUN": "3", "märkligt|ADV": "3", "uppehållstillstånd|NOUN": "3", "original|NOUN": "3", "utdelning|NOUN": "3", "julklapp|NOUN": "3", "klapp|NOUN": "3", "långvarig|ADJ": "3", "still|ADV": "3", "sammansättning|NOUN": "3", "oändlig|ADJ": "3", "oerhörd|ADJ": "3", "rast|NOUN": "3", "skapare|NOUN": "3", "benämning|NOUN": "3", "transportera|VERB": "3", "uppdelning|NOUN": "3", "väsen|NOUN": "3", "islamist|NOUN": "3", "självklarhet|NOUN": "3", "beaktande|NOUN": "3", "i kombination med|ADP": "3", "reta|VERB": "3", "trakt|NOUN": "3", "inledningsvis|ADV": "3", "krog|NOUN": "3", "enig|ADJ": "3", "ärva|VERB": "3", "jätte|NOUN": "3", "börda|NOUN": "3", "föregå|VERB": "3", "publicering|NOUN": "3", "skifte|NOUN": "3", "aktivist|NOUN": "3", "guide|NOUN": "3", "smälta|VERB": "3", "styrka|VERB": "3", "frysa|VERB": "3", "noggrann|ADJ": "3", "systematisk|ADJ": "3", "tillträde|NOUN": "3", "oväntat|ADV": "3", "kompetent|ADJ": "3", "prostitution|NOUN": "3", "skick|NOUN": "3", "mätt|ADJ": "3", "inköp|NOUN": "3", "ficka|NOUN": "3", "nederlag|NOUN": "3", "ansökning|NOUN": "3", "verkligt|ADV": "3", "story|NOUN": "3", "byrå|NOUN": "3", "dryck|NOUN": "3", "smidig|ADJ": "3", "synvinkel|NOUN": "3", "så gott som|ADV": "3", "försvaga|VERB": "3", "gräs|NOUN": "3", "förfluten|ADJ": "3", "simma|VERB": "3", "fysik|NOUN": "3", "hockey|NOUN": "3", "produktivitet|NOUN": "3", "incitament|NOUN": "3", "kontrast|NOUN": "3", "läpp|NOUN": "3", "progressiv|ADJ": "3", "anmärkningsvärd|ADJ": "3", "mobil|NOUN": "3", "tull|NOUN": "3", "fotografera (vardagl. fota)|VERB": "3", "skärm|NOUN": "3", "databas|NOUN": "3", "fynd|NOUN": "3", "bekymmer|NOUN": "3", "underhåll|NOUN": "3", "i gång (el. igång)|ADV": "3", "tätt|ADV": "3", "överlägsen|ADJ": "3", "grek|NOUN": "3", "kedja|NOUN": "3", "sår|NOUN": "3", "uppenbarelse|NOUN": "3", "utfall|NOUN": "3", "naiv|ADJ": "3", "still|ADJ": "3", "morgondag|NOUN": "3", "nöd|NOUN": "3", "motorväg|NOUN": "3", "utvecklingsland|NOUN": "3", "avhandling|NOUN": "3", "godis|NOUN": "3", "ko|NOUN": "3", "påvisa|VERB": "3", "trampa|VERB": "3", "ambassadör|NOUN": "3", "torka|VERB": "3", "så att säga|ADV": "3", "titt|NOUN": "3", "spränga|VERB": "3", "halva|NOUN": "3", "känneteckna|VERB": "3", "ombud|NOUN": "3", "ortodox|ADJ": "3", "problematisk|ADJ": "3", "virus|NOUN": "3", "himmelsk|ADJ": "3", "uppsats|NOUN": "3", "strålande|ADJ": "3", "bindande|ADJ": "3", "alltjämt|ADV": "3", "jämt|ADV": "3", "hungrig|ADJ": "3", "elak|ADJ": "3", "bosättning|NOUN": "3", "miljövänlig|ADJ": "3", "förfogande|NOUN": "3", "lucka|NOUN": "3", "procentenhet|NOUN": "3", "sammanträde|NOUN": "3", "musikalisk|ADJ": "3", "självförtroende|NOUN": "3", "cool|ADJ": "3", "fördjupa|VERB": "3", "ingång|NOUN": "3", "sed|NOUN": "3", "taxi|NOUN": "3", "vänja|VERB": "3", "författning|NOUN": "3", "huvudperson|NOUN": "3", "hypotes|NOUN": "3", "panik|NOUN": "3", "stämma|NOUN": "3", "avslutning|NOUN": "3", "deklaration|NOUN": "3", "sväng|NOUN": "3", "presidentval|NOUN": "3", "undgå|VERB": "3", "illusion|NOUN": "3", "international|NOUN": "3", "intrång|NOUN": "3", "skattepengar|NOUN": "3", "stolthet|NOUN": "3", "utnyttjande|NOUN": "3", "överlevnad|NOUN": "3", "problematik|NOUN": "3", "sällsynt|ADJ": "3", "dumhet|NOUN": "3", "flöde|NOUN": "3", "jättebra|ADJ": "3", "i jämförelse med|ADP": "3", "medborgarskap|NOUN": "3", "snack|NOUN": "3", "parallellt|ADV": "3", "påföljd|NOUN": "3", "söder om|ADP": "3", "strax efter|ADV": "3", "talang|NOUN": "3", "varmt|ADV": "3", "pjäs|NOUN": "3", "kansli|NOUN": "3", "lagligt|ADV": "3", "sand|NOUN": "3", "fildelare|NOUN": "3", "liga|NOUN": "3", "parlamentarisk|ADJ": "3", "vittnesbörd|NOUN": "3", "avrätta|VERB": "3", "fiske|NOUN": "3", "gynnsam|ADJ": "3", "dokumentär|NOUN": "3", "dödlig|ADJ": "3", "beteckning|NOUN": "3", "jämte|ADP": "3", "uttryckligen|ADV": "3", "distrikt|NOUN": "3", "påse|NOUN": "3", "baksida|NOUN": "3", "plånbok|NOUN": "3", "uppsägning|NOUN": "3", "fullfölja|VERB": "3", "foga|VERB": "3", "psykologi|NOUN": "3", "hjul|NOUN": "3", "klänning|NOUN": "3", "anteckning|NOUN": "3", "trä|NOUN": "3", "belägg|NOUN": "3", "blunda|VERB": "3", "vik|NOUN": "3", "bråk|NOUN": "3", "värva|VERB": "3", "biblisk|ADJ": "3", "sikta|VERB": "3", "uteslutande|ADV": "3", "pryl|NOUN": "3", "begravning|NOUN": "3", "naturligt|ADV": "3", "bredd|NOUN": "3", "frälsning|NOUN": "3", "funktionshinder|NOUN": "3", "såvida|SCONJ": "3", "avvika|VERB": "3", "influensa|NOUN": "3", "medvetenhet|NOUN": "3", "muskel|NOUN": "3", "ointressant|ADJ": "3", "samhällelig|ADJ": "3", "apropå|ADP": "3", "cirkel|NOUN": "3", "rekord|NOUN": "3", "bemärkelse|NOUN": "3", "djävul|NOUN": "3", "tålamod|NOUN": "3", "utspel|NOUN": "3", "verkställa|VERB": "3", "hjälpmedel|NOUN": "3", "riksdagsval|NOUN": "3", "svära|VERB": "3", "tagg|NOUN": "3", "deklarera|VERB": "3", "meningsfull|ADJ": "3", "i anslutning till|ADP": "3", "rimligen|ADV": "3", "minut (förk. min.)|NOUN": "3", "annanstans|ADV": "3", "knapp|ADJ": "3", "kvartal|NOUN": "3", "party|NOUN": "3", "imponera|VERB": "3", "innanför|ADP": "3", "expansion|NOUN": "3", "vaken|ADJ": "3", "kunnig|ADJ": "3", "scenario|NOUN": "3", "leverans|NOUN": "3", "medelstor|ADJ": "3", "salt|NOUN": "3", "sannolik|ADJ": "3", "vänskap|NOUN": "3", "farmor|NOUN": "3", "tiotusentals|ADV": "3", "lokalt|ADV": "3", "frigöra|VERB": "3", "prestation|NOUN": "3", "olämplig|ADJ": "3", "belöning|NOUN": "3", "styrning|NOUN": "3", "säte|NOUN": "3", "sjukförsäkring|NOUN": "3", "upplysa|VERB": "3", "halvtimme|NOUN": "3", "uppsättning|NOUN": "3", "sms|NOUN": "3", "elektrisk|ADJ": "3", "folkbildning|NOUN": "3", "kriminalitet|NOUN": "3", "födelse|NOUN": "3", "registrering|NOUN": "3", "nord|NOUN": "3", "färdas|VERB": "3", "världsbild|NOUN": "3", "brista|VERB": "3", "prinsessa|NOUN": "3", "överlåta|VERB": "3", "konsumera|VERB": "3", "vardaglig|ADJ": "3", "besättning|NOUN": "3", "manus|NOUN": "3", "mestadels|ADV": "3", "glädjande|ADJ": "3", "imperialism|NOUN": "3", "departement|NOUN": "3", "förfölja|VERB": "3", "operativ|ADJ": "3", "fullmäktige|NOUN": "3", "kommunfullmäktige|NOUN": "3", "nyliberal|ADJ": "3", "sparande|NOUN": "3", "interpellation|NOUN": "3", "marxism|NOUN": "3", "trång|ADJ": "3", "angelägenhet|NOUN": "3", "potatis|NOUN": "3", "medeltida|ADJ": "3", "underhållande|ADJ": "3", "ensamhet|NOUN": "3", "noggrant|ADV": "3", "sprit|NOUN": "3", "panna|NOUN": "3", "sakfråga|NOUN": "3", "brun|ADJ": "3", "kind|NOUN": "3", "förekomst|NOUN": "3", "härifrån|ADV": "3", "okunnig|ADJ": "3", "oförändrad|ADJ": "3", "sedermera|ADV": "3", "möjligtvis|ADV": "3", "fordra|VERB": "3", "förhållningssätt|NOUN": "3", "hall|NOUN": "3", "regelbunden|ADJ": "3", "klassiker|NOUN": "3", "uppkomst|NOUN": "3", "vägledning|NOUN": "3", "kika|VERB": "3", "dos|NOUN": "3", "försiktigt|ADV": "3", "blodig|ADJ": "3", "dynamisk|ADJ": "3", "portion|NOUN": "3", "smutsig|ADJ": "3", "svika|VERB": "3", "smått|ADV": "3", "bortsett från|ADP": "3", "förstärkning|NOUN": "3", "förteckning|NOUN": "3", "narkotikum|NOUN": "3", "björn|NOUN": "3", "engelsman|NOUN": "3", "utropa|VERB": "3", "fascism|NOUN": "3", "gnälla|VERB": "3", "underbart|ADV": "3", "ankomst|NOUN": "3", "barnbarn|NOUN": "3", "gudstjänst|NOUN": "3", "pott|NOUN": "3", "regissör|NOUN": "3", "turk|NOUN": "3", "hylla|NOUN": "3", "tillfälligt|ADV": "3", "ungdomsförbund|NOUN": "3", "eftersträva|VERB": "3", "förflytta|VERB": "3", "sekreterare|NOUN": "3", "missnöjd|ADJ": "3", "värdelös|ADJ": "3", "doft|NOUN": "3", "passiv|ADJ": "3", "uppfinning|NOUN": "3", "språklig|ADJ": "3", "härska|VERB": "3", "kast|NOUN": "3", "sympati|NOUN": "3", "behörighet|NOUN": "3", "förknippa|VERB": "3", "insändare|NOUN": "3", "judendom|NOUN": "3", "sjuksköterska|NOUN": "3", "tält|NOUN": "3", "uppgång|NOUN": "3", "inskränka|VERB": "3", "prestera|VERB": "3", "udda|ADJ": "3", "journal|NOUN": "3", "diplomatisk|ADJ": "3", "tillfredsställande|ADJ": "3", "förakt|NOUN": "3", "regera|VERB": "3", "indirekt|ADJ": "3", "gyllene|ADJ": "3", "söderut|ADV": "3", "kapitalist|NOUN": "3", "genomslag|NOUN": "3", "teologisk|ADJ": "3", "matta|NOUN": "3", "medelklass|NOUN": "3", "målgrupp|NOUN": "3", "sortera|VERB": "3", "säkerhetspolitik|NOUN": "3", "födelsedag|NOUN": "3", "misshandla|VERB": "3", "mynt|NOUN": "3", "rörlig|ADJ": "3", "gods|NOUN": "3", "beredning|NOUN": "3", "traditionellt|ADV": "3", "bliva|VERB": "3", "agent|NOUN": "3", "exklusiv|ADJ": "3", "handlande|NOUN": "3", "socker|NOUN": "3", "upplopp|NOUN": "3", "kaka|NOUN": "3", "kollektivtrafik|NOUN": "3", "anlägga|VERB": "3", "upphandling|NOUN": "3", "breda|VERB": "3", "realitet|NOUN": "4", "marknadsföra|VERB": "4", "vitt|ADV": "4", "vrede|NOUN": "4", "satan|NOUN": "4", "statistisk|ADJ": "4", "ödmjuk|ADJ": "4", "i natt|ADV": "4", "klarhet|NOUN": "4", "långsiktigt|ADV": "4", "anstränga|VERB": "4", "generös|ADJ": "4", "mellanrum|NOUN": "4", "sken|NOUN": "4", "upplösning|NOUN": "4", "vistelse|NOUN": "4", "växla|VERB": "4", "strukturell|ADJ": "4", "förvärva|VERB": "4", "regi|NOUN": "4", "anka|NOUN": "4", "redogörelse|NOUN": "4", "statsmakt|NOUN": "4", "etta|NOUN": "4", "relativ|ADJ": "4", "vindkraft|NOUN": "4", "imperialistisk|ADJ": "4", "måltid|NOUN": "4", "till synes|ADV": "4", "belöna|VERB": "4", "importera|VERB": "4", "liter|NOUN": "4", "rentav|ADV": "4", "stormakt|NOUN": "4", "samtida|ADJ": "4", "legal|ADJ": "4", "principiell|ADJ": "4", "valfrihet|NOUN": "4", "tydlighet|NOUN": "4", "växthusgas|NOUN": "4", "evenemang|NOUN": "4", "lösenord|NOUN": "4", "dialekt|NOUN": "4", "behärska|VERB": "4", "föregångare|NOUN": "4", "homosexualitet|NOUN": "4", "seg|ADJ": "4", "licens|NOUN": "4", "platt|ADJ": "4", "iver|NOUN": "4", "resenär|NOUN": "4", "utrota|VERB": "4", "uppfinna|VERB": "4", "cup|NOUN": "4", "omvänd|ADJ": "4", "dagordning|NOUN": "4", "perfekt|ADV": "4", "splittring|NOUN": "4", "inbilla|VERB": "4", "avge|VERB": "4", "partnerskap|NOUN": "4", "löna sig|VERB": "4", "brutal|ADJ": "4", "konstruera|VERB": "4", "ärlighet|NOUN": "4", "bekväm|ADJ": "4", "presskonferens|NOUN": "4", "osannolik|ADJ": "4", "totalitär|ADJ": "4", "åtgärda|VERB": "4", "flickvän|NOUN": "4", "norrut|ADV": "4", "arbetstillfälle|NOUN": "4", "inträde|NOUN": "4", "släpa|VERB": "4", "övervägande|NOUN": "4", "skilsmässa|NOUN": "4", "utforska|VERB": "4", "bildande|ADJ": "4", "tyngd|NOUN": "4", "frälsare|NOUN": "4", "invadera|VERB": "4", "personuppgift|NOUN": "4", "förhand|NOUN": "4", "gruppering|NOUN": "4", "tekniskt|ADV": "4", "dagstidning|NOUN": "4", "oacceptabel|ADJ": "4", "serb|NOUN": "4", "flytande|ADJ": "4", "justera|VERB": "4", "adel|NOUN": "4", "konsult|NOUN": "4", "nervös|ADJ": "4", "sekt|NOUN": "4", "slöja|NOUN": "4", "välkommen|INTJ": "4", "läcka|VERB": "4", "afton|NOUN": "4", "introduktion|NOUN": "4", "livstid|NOUN": "4", "demonstrant|NOUN": "4", "flexibilitet|NOUN": "4", "hed|NOUN": "4", "kol|NOUN": "4", "uppväxt|NOUN": "4", "efterlysa|VERB": "4", "grönsak|NOUN": "4", "samordna|VERB": "4", "järn|NOUN": "4", "distribution|NOUN": "4", "automatisk|ADJ": "4", "transaktion|NOUN": "4", "däck|NOUN": "4", "observation|NOUN": "4", "typiskt|ADV": "4", "inskränkning|NOUN": "4", "mata|VERB": "4", "paradis|NOUN": "4", "ingenjör|NOUN": "4", "koncentration|NOUN": "4", "plus|NOUN": "4", "dugg|NOUN": "4", "samtid|NOUN": "4", "uppståndelse|NOUN": "4", "slaveri|NOUN": "4", "ålägga|VERB": "4", "framkalla|VERB": "4", "utkast|NOUN": "4", "framträdande|ADJ": "4", "desperat|ADJ": "4", "någon som helst|DET": "4", "flitigt|ADV": "4", "offensiv|NOUN": "4", "sångare|NOUN": "4", "ingrepp|NOUN": "4", "otalig|ADJ": "4", "diagram|NOUN": "4", "inbjuda|VERB": "4", "motivation|NOUN": "4", "utplåna|VERB": "4", "gymnasieskola|NOUN": "4", "bearbeta|VERB": "4", "förlåtelse|NOUN": "4", "snurra|VERB": "4", "skildring|NOUN": "4", "sändning|NOUN": "4", "baby|NOUN": "4", "förvara|VERB": "4", "rabatt|NOUN": "4", "rota|VERB": "4", "apa|NOUN": "4", "sammanställa|VERB": "4", "stirra|VERB": "4", "avgörande|NOUN": "4", "manifestation|NOUN": "4", "uppenbara|VERB": "4", "maila|VERB": "4", "medmänniska|NOUN": "4", "genombrott|NOUN": "4", "proletär|ADJ": "4", "fika|NOUN": "4", "spaning|NOUN": "4", "beordra|VERB": "4", "förbinda|VERB": "4", "jämförbar|ADJ": "4", "socialt|ADV": "4", "fullgöra|VERB": "4", "förr eller senare|ADV": "4", "palm|NOUN": "4", "förvirring|NOUN": "4", "privatisering|NOUN": "4", "chock|NOUN": "4", "oundviklig|ADJ": "4", "samtycke|NOUN": "4", "förband|NOUN": "4", "missbruka|VERB": "4", "förvärra|VERB": "4", "investerare|NOUN": "4", "vackert|ADV": "4", "utbredd|ADJ": "4", "bio|NOUN": "4", "oförmåga|NOUN": "4", "sammanlagd|ADJ": "4", "klippa|NOUN": "4", "cd|NOUN": "4", "knut|NOUN": "4", "fras|NOUN": "4", "indikera|VERB": "4", "vardera|PRON": "4", "arrangör|NOUN": "4", "profetia|NOUN": "4", "därutöver|ADV": "4", "förnya|VERB": "4", "hederlig|ADJ": "4", "inhämta|VERB": "4", "skånsk|ADJ": "4", "abstrakt|ADJ": "4", "dämpa|VERB": "4", "tillhörighet|NOUN": "4", "möbel|NOUN": "4", "ringa|ADJ": "4", "sky|NOUN": "4", "anvisning|NOUN": "4", "hatt|NOUN": "4", "tokig|ADJ": "4", "förvärv|NOUN": "4", "med flera (förk. m.fl., m fl)|ADV": "4", "omgående|ADV": "4", "bedrägeri|NOUN": "4", "mobilisera|VERB": "4", "signatur|NOUN": "4", "skälig|ADJ": "4", "expandera|VERB": "4", "förkunna|VERB": "4", "böja|VERB": "4", "förenkla|VERB": "4", "viga|VERB": "4", "justitieminister|NOUN": "4", "fjärdedel|NOUN": "4", "substans|NOUN": "4", "tömma|VERB": "4", "utmärka|VERB": "4", "ende|ADJ": "4", "förnyelse|NOUN": "4", "subjektiv|ADJ": "4", "burk|NOUN": "4", "human|ADJ": "4", "mista|VERB": "4", "sanktion|NOUN": "4", "fler och fler|PRON": "4", "omsättning|NOUN": "4", "besitta|VERB": "4", "initiera|VERB": "4", "skrivande|NOUN": "4", "hänseende|NOUN": "4", "härstamma|VERB": "4", "censur|NOUN": "4", "kollektiv|NOUN": "4", "promenera|VERB": "4", "supa|VERB": "4", "legitimitet|NOUN": "4", "befäl|NOUN": "4", "sökande|NOUN": "4", "pojkvän|NOUN": "4", "poängtera|VERB": "4", "överträdelse|NOUN": "4", "klimatfråga|NOUN": "4", "telefonsamtal|NOUN": "4", "beredskap|NOUN": "4", "vers|NOUN": "4", "monarki|NOUN": "4", "ockupera|VERB": "4", "skum|ADJ": "4", "turism|NOUN": "4", "befrielse|NOUN": "4", "byxa|NOUN": "4", "rekrytera|VERB": "4", "förmögenhet|NOUN": "4", "gången|ADJ": "4", "liksom|SCONJ": "4", "äpple|NOUN": "4", "höjdpunkt|NOUN": "4", "sammanställning|NOUN": "4", "underhållning|NOUN": "4", "uppbyggnad|NOUN": "4", "etablissemang|NOUN": "4", "kontinuerligt|ADV": "4", "krama|VERB": "4", "missförstånd|NOUN": "4", "nationalistisk|ADJ": "4", "obalans|NOUN": "4", "nyår|NOUN": "4", "produktiv|ADJ": "4", "till rätta|ADV": "4", "avveckling|NOUN": "4", "provocera|VERB": "4", "erfaren|ADJ": "4", "blank|ADJ": "4", "singel|NOUN": "4", "försörjning|NOUN": "4", "irländsk|ADJ": "4", "kurd|NOUN": "4", "psykolog|NOUN": "4", "samtala|VERB": "4", "sekel|NOUN": "4", "federal|ADJ": "4", "frustration|NOUN": "4", "fundamental|ADJ": "4", "omge|VERB": "4", "företa|VERB": "4", "utdrag|NOUN": "4", "fram och tillbaka|ADV": "4", "lågt|ADV": "4", "skal|NOUN": "4", "irakisk|ADJ": "4", "parallell|NOUN": "4", "avslag|NOUN": "4", "emellanåt|ADV": "4", "källare|NOUN": "4", "merpart|NOUN": "4", "vetskap|NOUN": "4", "delägare|NOUN": "4", "distans|NOUN": "4", "eliminera|VERB": "4", "i motsats till|ADP": "4", "tolerans|NOUN": "4", "krigare|NOUN": "4", "bosätta|VERB": "4", "filma|VERB": "4", "upplägg|NOUN": "4", "föda|NOUN": "4", "överläggning|NOUN": "4", "miss|NOUN": "4", "moské|NOUN": "4", "passion|NOUN": "4", "zon|NOUN": "4", "tunga|NOUN": "4", "vass|ADJ": "4", "klient|NOUN": "4", "spana|VERB": "4", "utbetalning|NOUN": "4", "obetydlig|ADJ": "4", "kurdisk|ADJ": "4", "relevans|NOUN": "4", "förutsatt att|SCONJ": "4", "motarbeta|VERB": "4", "påtryckning|NOUN": "4", "efterföljande|ADJ": "4", "nyhetsbrev|NOUN": "4", "årsskifte|NOUN": "4", "avvikelse|NOUN": "4", "tilltala|VERB": "4", "stift|NOUN": "4", "hemlös|ADJ": "4", "splittra|VERB": "4", "bosätta sig|VERB": "4", "bekräftelse|NOUN": "4", "försvarsminister|NOUN": "4", "dokumentera|VERB": "4", "lydnad|NOUN": "4", "tragedi|NOUN": "4", "organism|NOUN": "4", "socialtjänst|NOUN": "4", "tillskriva|VERB": "4", "humanist|NOUN": "4", "snett|ADV": "4", "firma|NOUN": "4", "förankring|NOUN": "4", "reporänta|NOUN": "4", "sekulär|ADJ": "4", "fortsättningsvis|ADV": "4", "erfara|VERB": "4", "inblandning|NOUN": "4", "signalspaning|NOUN": "4", "svininfluensa|NOUN": "4", "liknelse|NOUN": "4", "beväpnad|ADJ": "4", "härligt|ADV": "4", "ingripande|NOUN": "4", "pigg|ADJ": "4", "bebyggelse|NOUN": "4", "fysiskt|ADV": "4", "romantisk|ADJ": "4", "ingående|ADJ": "4", "märkning|NOUN": "4", "lojalitet|NOUN": "4", "penna|NOUN": "4", "får|NOUN": "4", "illustration|NOUN": "4", "rock|NOUN": "4", "innehav|NOUN": "4", "tilltro|NOUN": "4", "dvd|NOUN": "4", "bensin|NOUN": "4", "bromsa|VERB": "4", "bråka|VERB": "4", "kula|NOUN": "4", "svält|NOUN": "4", "klo|NOUN": "4", "sektion|NOUN": "4", "avskaffande|NOUN": "4", "examen|NOUN": "4", "religionsfrihet|NOUN": "4", "utåt|ADV": "4", "balansera|VERB": "4", "heltid|NOUN": "4", "hemifrån|ADV": "4", "stifta|VERB": "4", "verkställande|ADJ": "4", "asyl|NOUN": "4", "graviditet|NOUN": "4", "korsa|VERB": "4", "avlägsna|VERB": "4", "beställning|NOUN": "4", "fasad|NOUN": "4", "infinna sig|VERB": "4", "hyfsat|ADV": "4", "julafton|NOUN": "4", "organisk|ADJ": "4", "åtnjuta|VERB": "4", "för alltid|ADV": "4", "hemmaplan|NOUN": "4", "kloster|NOUN": "4", "förlita sig|VERB": "4", "förlägga|VERB": "4", "spontan|ADJ": "4", "informell|ADJ": "4", "förvåning|NOUN": "4", "iaktta|VERB": "4", "körkort|NOUN": "4", "försäkringsbolag|NOUN": "4", "missnöje|NOUN": "4", "etnicitet|NOUN": "4", "inbjudan|NOUN": "4", "dyster|ADJ": "4", "okunskap|NOUN": "4", "garanterat|ADV": "4", "sammanfattningsvis|ADV": "4", "spark|NOUN": "4", "arbetsdag|NOUN": "4", "silver|NOUN": "4", "organisatorisk|ADJ": "4", "slutgiltig|ADJ": "4", "tungt|ADV": "4", "bekänna|VERB": "4", "kostym|NOUN": "4", "schema|NOUN": "4", "långtgående|ADJ": "4", "mask|NOUN": "4", "materiel|NOUN": "4", "mobbning|NOUN": "4", "leksak|NOUN": "4", "spridd|ADJ": "4", "stava|VERB": "4", "tillit|NOUN": "4", "modig|ADJ": "4", "utbrott|NOUN": "4", "apparat|NOUN": "4", "disk|NOUN": "4", "drama|NOUN": "4", "exportera|VERB": "4", "försoning|NOUN": "4", "universell|ADJ": "4", "beroende|NOUN": "4", "surfa|VERB": "4", "diktator|NOUN": "4", "passage|NOUN": "4", "inbyggd|ADJ": "4", "plåga|VERB": "4", "strikt|ADJ": "4", "utlova|VERB": "4", "riksbank|NOUN": "4", "återta|VERB": "4", "dokumentation|NOUN": "4", "ingrediens|NOUN": "4", "inträda|VERB": "4", "show|NOUN": "4", "bak|ADV": "4", "delaktighet|NOUN": "4", "i viss mån|ADV": "4", "odling|NOUN": "4", "vardagsrum|NOUN": "4", "fascinerande|ADJ": "4", "kontext|NOUN": "4", "lina|NOUN": "4", "folkhögskola|NOUN": "4", "glasögon|NOUN": "4", "inviga|VERB": "4", "rop|NOUN": "4", "varannan|DET": "4", "disciplin|NOUN": "4", "europé|NOUN": "4", "härskare|NOUN": "4", "återkomst|NOUN": "4", "i fred|ADV": "4", "kompensation|NOUN": "4", "representativ|ADJ": "4", "strömma|VERB": "4", "kartlägga|VERB": "4", "systematiskt|ADV": "4", "i relation till|ADP": "4", "uppe|PART": "4", "yxa|NOUN": "4", "bevakning|NOUN": "4", "missionär|NOUN": "4", "rätta|NOUN": "4", "bekännelse|NOUN": "4", "ensidig|ADJ": "4", "högtid|NOUN": "4", "institutionell|ADJ": "4", "psykiskt|ADV": "4", "skjorta|NOUN": "4", "under förutsättning att|SCONJ": "4", "rehabilitering|NOUN": "4", "skärgård|NOUN": "4", "övervinna|VERB": "4", "enkät|NOUN": "4", "garderob|NOUN": "4", "läxa|NOUN": "4", "med avseende på|ADP": "4", "trumma|NOUN": "4", "pol|NOUN": "4", "choklad|NOUN": "4", "återhämtning|NOUN": "4", "bakterie|NOUN": "4", "exploatering|NOUN": "4", "kärnkraftverk|NOUN": "4", "stig|NOUN": "4", "primär|ADJ": "4", "republikan|NOUN": "4", "gestalt|NOUN": "4", "konstitutionell|ADJ": "4", "avslutningsvis|ADV": "4", "indian|NOUN": "4", "ingenstans|ADV": "4", "nuförtiden (el. nu för tiden)|ADV": "4", "runda|NOUN": "4", "baltisk|ADJ": "4", "farfar|NOUN": "4", "förtydliga|VERB": "4", "gärningsman|NOUN": "4", "succé|NOUN": "4", "tröst|NOUN": "4", "epok|NOUN": "4", "intention|NOUN": "4", "nedskärning|NOUN": "4", "tillika|ADV": "4", "remiss|NOUN": "4", "skåda|VERB": "4", "bevittna|VERB": "4", "främling|NOUN": "4", "juridik|NOUN": "4", "utvisning|NOUN": "4", "folkrätt|NOUN": "4", "legitim|ADJ": "4", "bostadsområde|NOUN": "4", "egyptisk|ADJ": "4", "glatt|ADV": "4", "hyresgäst|NOUN": "4", "radikalt|ADV": "4", "vinge|NOUN": "4", "klassa|VERB": "4", "legend|NOUN": "4", "öre|NOUN": "4", "nazistisk|ADJ": "4", "varsin|PRON": "4", "begrava|VERB": "4", "funktionsnedsättning|NOUN": "4", "kontra|ADP": "4", "persisk|ADJ": "4", "tillskott|NOUN": "4", "klagomål|NOUN": "4", "konstverk|NOUN": "4", "kortsiktig|ADJ": "4", "avliden|ADJ": "6", "backe|NOUN": "4", "förespråkare|NOUN": "4", "indikator|NOUN": "4", "nutida|ADJ": "4", "textstorlek|NOUN": "4", "åta|VERB": "4", "asiatisk|ADJ": "4", "meny|NOUN": "4", "muntlig|ADJ": "4", "nedre|ADJ": "4", "regeringsform|NOUN": "4", "otrevlig|ADJ": "4", "publikation|NOUN": "4", "halt|NOUN": "4", "borg|NOUN": "4", "pedofil|NOUN": "4", "porträtt|NOUN": "4", "utomstående|ADJ": "4", "ironi|NOUN": "4", "manipulera|VERB": "4", "afghansk|ADJ": "4", "jag|NOUN": "4", "utomhus|ADV": "4", "privilegium|NOUN": "4", "rensning|NOUN": "4", "etapp|NOUN": "4", "minimera|VERB": "4", "till fullo|ADV": "4", "representation|NOUN": "4", "latin|NOUN": "4", "måhända|ADV": "4", "serbisk|ADJ": "4", "estetisk|ADJ": "4", "explodera|VERB": "4", "folkrörelse|NOUN": "4", "grundare|NOUN": "4", "konspiration|NOUN": "4", "kritiskt|ADV": "4", "kurva|NOUN": "4", "operera|VERB": "4", "turné|NOUN": "4", "åskådare|NOUN": "4", "forntid|NOUN": "4", "alliansregering|NOUN": "4", "framgångsrikt|ADV": "4", "ovan|ADP": "4", "robot|NOUN": "4", "försvarare|NOUN": "4", "landslag|NOUN": "4", "proportion|NOUN": "4", "verkstad|NOUN": "4", "ask|NOUN": "4", "bomba|VERB": "4", "jeans|NOUN": "4", "jordbävning|NOUN": "4", "ratt|NOUN": "4", "brant|ADJ": "4", "befälhavare|NOUN": "4", "bot|NOUN": "4", "dusch|NOUN": "4", "konsensus|NOUN": "4", "könsneutral|ADJ": "4", "våldta|VERB": "4", "skruva|VERB": "4", "slutföra|VERB": "4", "återspegla|VERB": "4", "eko|NOUN": "4", "horisont|NOUN": "4", "inkomma|VERB": "4", "ministerråd|NOUN": "4", "beslutsfattare|NOUN": "4", "suck|NOUN": "4", "utlösa|VERB": "4", "flygbolag|NOUN": "4", "spegel|NOUN": "4", "konventionell|ADJ": "4", "metall|NOUN": "4", "återstående|ADJ": "4", "i fjol|ADV": "4", "lönsamhet|NOUN": "4", "vari|ADV": "4", "balanserad|ADJ": "4", "antiken|NOUN": "4", "innovativ|ADJ": "4", "utnämna|VERB": "4", "islamistisk|ADJ": "4", "pricka|VERB": "4", "tunnel|NOUN": "4", "avreglering|NOUN": "4", "bristfällig|ADJ": "4", "ensamstående|ADJ": "4", "inomhus|ADV": "4", "kapabel|ADJ": "4", "autonom|ADJ": "4", "mekanisk|ADJ": "4", "övertygande|ADJ": "4", "kvarvarande|ADJ": "4", "vägnar|NOUN": "4", "befara|VERB": "4", "beundra|VERB": "4", "förfall|NOUN": "4", "toppmöte|NOUN": "4", "trakasseri|NOUN": "4", "kupp|NOUN": "4", "bistå|VERB": "4", "sno|VERB": "4", "genuin|ADJ": "4", "nuläge|NOUN": "4", "ros|NOUN": "4", "tittare|NOUN": "4", "trasig|ADJ": "4", "check|NOUN": "4", "irrelevant|ADJ": "4", "moraliskt|ADV": "4", "överlag|ADV": "4", "förstånd|NOUN": "4", "blockad|NOUN": "4", "nutid|NOUN": "4", "omställning|NOUN": "4", "rumpa|NOUN": "4", "förebyggande|ADJ": "4", "notis|NOUN": "4", "mejl|NOUN": "4", "moms|NOUN": "4", "samspel|NOUN": "4", "aktiebolag|NOUN": "4", "jävel|NOUN": "4", "ledighet|NOUN": "4", "prat|NOUN": "4", "uppför|ADP": "4", "riksdagsbeslut|NOUN": "4", "balkong|NOUN": "4", "glass|NOUN": "4", "kallelse|NOUN": "4", "omsätta|VERB": "4", "destruktiv|ADJ": "4", "för|NOUN": "4", "sy|VERB": "4", "virtuell|ADJ": "4", "ärkebiskop|NOUN": "4", "invända|VERB": "4", "restriktion|NOUN": "4", "snar|ADJ": "4", "upprörd|ADJ": "4", "koncern|NOUN": "4", "minimal|ADJ": "4", "konvent|NOUN": "4", "fientlig|ADJ": "4", "förfader|NOUN": "4", "underhålla|VERB": "4", "vansinnig|ADJ": "4", "biografi|NOUN": "4", "räddning|NOUN": "4", "rör|NOUN": "4", "fiska|VERB": "4", "försämring|NOUN": "4", "mode|NOUN": "4", "programledare|NOUN": "4", "ytlig|ADJ": "4", "genomgående|ADJ": "4", "tron|NOUN": "4", "efternamn|NOUN": "4", "hämnd|NOUN": "4", "puls|NOUN": "4", "tidsperiod|NOUN": "4", "medelålder|NOUN": "4", "nyfikenhet|NOUN": "4", "barnomsorg|NOUN": "4", "ggr (gånger)|NOUN": "4", "framstående|ADJ": "4", "innehavare|NOUN": "4", "funktionshindrad|ADJ": "4", "isolering|NOUN": "4", "kreditkort|NOUN": "4", "otillräcklig|ADJ": "4", "arbetsmiljö|NOUN": "4", "fusk|NOUN": "4", "lik|NOUN": "4", "nationalitet|NOUN": "4", "smör|NOUN": "4", "tillträda|VERB": "4", "bänk|NOUN": "4", "korthet|NOUN": "4", "kungarike|NOUN": "4", "målvakt|NOUN": "4", "svans|NOUN": "4", "utvisa|VERB": "4", "lite grann|ADV": "4", "efterträdare|NOUN": "4", "närstående|ADJ": "4", "parallell|ADJ": "4", "plötslig|ADJ": "4", "rök|NOUN": "4", "skälla|VERB": "4", "valp|NOUN": "4", "fruktan|NOUN": "4", "rekrytering|NOUN": "4", "förövare|NOUN": "4", "popularitet|NOUN": "4", "symbolisera|VERB": "4", "kollaps|NOUN": "4", "kändis|NOUN": "4", "ont|NOUN": "4", "termin|NOUN": "4", "tills vidare|ADV": "4", "dilemma|NOUN": "4", "smärtsam|ADJ": "4", "holländsk|ADJ": "4", "klämma|VERB": "4", "ateist|NOUN": "4", "fotnot|NOUN": "4", "samverka|VERB": "4", "antik|ADJ": "4", "krånglig|ADJ": "4", "förpackning|NOUN": "4", "överskrida|VERB": "4", "aktivera|VERB": "4", "flytt|NOUN": "4", "vida|ADV": "4", "älg|NOUN": "4", "förstörelse|NOUN": "4", "elegant|ADJ": "4", "avgång|NOUN": "4", "montera|VERB": "4", "polisman|NOUN": "4", "preliminär|ADJ": "4", "primitiv|ADJ": "4", "avrättning|NOUN": "4", "nedåt|ADV": "4", "real|ADJ": "4", "överväldigande|ADJ": "4", "gym|NOUN": "4", "federation|NOUN": "4", "mötesplats|NOUN": "4", "öster|NOUN": "4", "beslutsfattande|NOUN": "4", "psykiatri|NOUN": "4", "handläggning|NOUN": "4", "utbryta|VERB": "4", "fientlighet|NOUN": "4", "inredning|NOUN": "4", "troll|NOUN": "4", "identisk|ADJ": "4", "riksförbund|NOUN": "4", "sal|NOUN": "4", "förtjust|ADV": "4", "generalsekreterare|NOUN": "4", "genomsyra|VERB": "4", "öppning|NOUN": "4", "obefintlig|ADJ": "4", "tillförlitlig|ADJ": "4", "näringsminister|NOUN": "4", "protein|NOUN": "4", "applåd|NOUN": "4", "ersättare|NOUN": "4", "onödigt|ADV": "4", "tjänstgöra|VERB": "4", "fastslå|VERB": "4", "slut|ADJ": "4", "solig|ADJ": "4", "gåta|NOUN": "4", "härlighet|NOUN": "4", "återuppta|VERB": "4", "fördriva|VERB": "4", "hertig|NOUN": "4", "påsk|NOUN": "4", "komplement|NOUN": "4", "modersmål|NOUN": "4", "beröm|NOUN": "4", "frö|NOUN": "4", "installation|NOUN": "4", "släcka|VERB": "4", "odds|NOUN": "4", "årsmöte|NOUN": "4", "arm|ADJ": "4", "kommunstyrelse|NOUN": "4", "mångkulturell|ADJ": "4", "varaktig|ADJ": "4", "horn|NOUN": "4", "sedel|NOUN": "4", "valsedel|NOUN": "4", "merit|NOUN": "4", "skinn|NOUN": "4", "badrum|NOUN": "4", "inbegripa|VERB": "4", "sovrum|NOUN": "4", "uppehålla|VERB": "4", "opassande|ADJ": "4", "hårddisk|NOUN": "4", "insamling|NOUN": "4", "oändligt|ADV": "4", "påminnelse|NOUN": "4", "marin|ADJ": "4", "opera|NOUN": "4", "aktieägare|NOUN": "4", "panel|NOUN": "4", "på något vis|ADV": "4", "inflytelserik|ADJ": "4", "polismyndighet|NOUN": "4", "vetenskapsman|NOUN": "4", "begåvad|ADJ": "4", "miljöfråga|NOUN": "4", "miste|PART": "4", "nicka|VERB": "4", "övervägande|ADJ": "4", "förtjänst|NOUN": "4", "inge|VERB": "4", "stolt|ADV": "4", "undergång|NOUN": "4", "ambitiös|ADJ": "4", "hebreisk|ADJ": "4", "växelkurs|NOUN": "4", "möda|NOUN": "4", "anklagad|ADJ": "4", "klassrum|NOUN": "4", "kontinuerlig|ADJ": "4", "si|ADV": "4", "entusiasm|NOUN": "4", "respons|NOUN": "4", "monster|NOUN": "4", "rån|NOUN": "4", "självkänsla|NOUN": "4", "sammanhållning|NOUN": "4", "sammanfalla|VERB": "4", "bara|SCONJ": "4", "intensivt|ADV": "4", "optimal|ADJ": "4", "suverän|ADJ": "4", "upp och ner|ADV": "4", "apotek|NOUN": "4", "hälla|VERB": "4", "käka|VERB": "4", "fäste|NOUN": "4", "hastigt|ADV": "4", "livslång|ADJ": "4", "svälta|VERB": "4", "välta|VERB": "4", "arbetsgivaravgift|NOUN": "4", "demon|NOUN": "4", "fastighetsskatt|NOUN": "4", "korridor|NOUN": "4", "stridsvagn|NOUN": "4", "tillvara|PART": "4", "vittnesmål|NOUN": "4", "ansvarsfull|ADJ": "4", "bagage|NOUN": "4", "evigt|ADV": "4", "koldioxidutsläpp|NOUN": "4", "fängsla|VERB": "4", "utflykt|NOUN": "4", "gratulera|VERB": "4", "studerande|NOUN": "4", "upprop|NOUN": "4", "utgåva|NOUN": "4", "vädja|VERB": "4", "finländsk|ADJ": "4", "morfar|NOUN": "4", "norrman|NOUN": "4", "skandinavisk|ADJ": "4", "tumme|NOUN": "4", "utslag|NOUN": "4", "familjemedlem|NOUN": "4", "lasta|VERB": "4", "ledarsida|NOUN": "4", "skräp|NOUN": "4", "smitta|VERB": "4", "påtala|VERB": "4", "stort|ADV": "4", "levnadsstandard|NOUN": "4", "palats|NOUN": "4", "tyska|NOUN": "4", "opinionsundersökning|NOUN": "4", "vetenskapligt|ADV": "4", "revidera|VERB": "4", "lovande|ADJ": "4", "orolighet|NOUN": "4", "brud|NOUN": "4", "tillvägagångssätt|NOUN": "4", "klistra|VERB": "4", "trams|NOUN": "4", "isär|PART": "4", "kärleksfull|ADJ": "4", "usch|INTJ": "4", "avslöjande|NOUN": "4", "beskatta|VERB": "4", "skrivbord|NOUN": "4", "utrikespolitisk|ADJ": "4", "vakta|VERB": "4", "arbetskamrat|NOUN": "4", "idiotisk|ADJ": "4", "spontant|ADV": "4", "tillställning|NOUN": "4", "tvärs|ADV": "4", "budgetår|NOUN": "4", "förtrycka|VERB": "4", "passande|ADJ": "4", "atom|NOUN": "4", "avta|VERB": "4", "chips|NOUN": "4", "markering|NOUN": "4", "tillåten|ADJ": "4", "öken|NOUN": "4", "sammanhängande|ADJ": "4", "fläck|NOUN": "4", "retorisk|ADJ": "4", "borgmästare|NOUN": "4", "förlorare|NOUN": "4", "melodi|NOUN": "4", "senat|NOUN": "4", "skarpt|ADV": "4", "sjöman|NOUN": "4", "bläddra|VERB": "4", "bärare|NOUN": "4", "gissning|NOUN": "4", "i onödan|ADV": "4", "stryk|NOUN": "4", "strålning|NOUN": "4", "terräng|NOUN": "4", "väva|VERB": "4", "skönt|ADV": "4", "spricka|VERB": "4", "äldreomsorg|NOUN": "4", "övertala|VERB": "4", "känslomässig|ADJ": "4", "feber|NOUN": "4", "härja|VERB": "4", "spelregel|NOUN": "4", "bekymrad|ADJ": "4", "annonsera|VERB": "4", "belastning|NOUN": "4", "flock|NOUN": "4", "inspektion|NOUN": "4", "laddning|NOUN": "4", "sammanslutning|NOUN": "4", "svek|NOUN": "4", "aska|NOUN": "4", "bekymra|VERB": "4", "finanspolitik|NOUN": "4", "godtycklig|ADJ": "4", "bluff|NOUN": "4", "distribuera|VERB": "4", "from|ADJ": "4", "förlopp|NOUN": "4", "nedläggning|NOUN": "4", "bestrida|VERB": "4", "huvudman|NOUN": "4", "ikapp|PART": "4", "empati|NOUN": "4", "sammansatt|ADJ": "4", "avlyssning|NOUN": "4", "dessförinnan|ADV": "4", "golf|NOUN": "4", "rasande|ADJ": "4", "reaktionär|ADJ": "4", "vifta|VERB": "4", "överklagande|NOUN": "4", "anor|NOUN": "4", "dominans|NOUN": "4", "lax|NOUN": "4", "organisering|NOUN": "4", "gift|NOUN": "4", "prostituerad|ADJ": "4", "återupprätta|VERB": "4", "hacka|VERB": "4", "medial|ADJ": "4", "entré|NOUN": "4", "farbror|NOUN": "4", "livlig|ADJ": "4", "packning|NOUN": "4", "essä|NOUN": "4", "magi|NOUN": "4", "självständigt|ADV": "4", "trötthet|NOUN": "4", "konsekvent|ADJ": "4", "rådgivning|NOUN": "4", "smälla|VERB": "4", "journalistisk|ADJ": "4", "officerare|NOUN": "4", "tjuv|NOUN": "4", "vidd|NOUN": "4", "belysning|NOUN": "4", "hänföra|VERB": "4", "nationalstat|NOUN": "4", "nedladdning|NOUN": "4", "växthuseffekt|NOUN": "4", "grotta|NOUN": "4", "matematisk|ADJ": "4", "ovanpå|ADP": "4", "pärla|NOUN": "4", "värk|NOUN": "4", "halvlek|NOUN": "4", "påtagligt|ADV": "4", "benägen|ADJ": "4", "recensera|VERB": "4", "diskriminera|VERB": "4", "pilot|NOUN": "4", "eftertanke|NOUN": "4", "fiktiv|ADJ": "4", "närliggande|ADJ": "4", "pålitlig|ADJ": "4", "korv|NOUN": "4", "reformera|VERB": "4", "pop|NOUN": "4", "fördubbla|VERB": "4", "militant|ADJ": "4", "sammantaget|ADV": "4", "tillkomst|NOUN": "4", "incident|NOUN": "4", "intill|ADV": "4", "underrättelse|NOUN": "4", "redigera|VERB": "4", "stadigt|ADV": "4", "baka|VERB": "4", "gud|INTJ": "4", "herregud|INTJ": "4", "observatör|NOUN": "4", "facit|NOUN": "4", "gruva|NOUN": "4", "obekväm|ADJ": "4", "fossil|ADJ": "4", "verkning|NOUN": "4", "kompromissa|VERB": "4", "konspirationsteori|NOUN": "4", "nacke|NOUN": "4", "svälja|VERB": "4", "tillstyrka|VERB": "4", "rättfärdighet|NOUN": "4", "adressat|NOUN": "4", "frågetecken|NOUN": "4", "image|NOUN": "4", "njutning|NOUN": "4", "utmärkt|ADV": "4", "isländsk|ADJ": "4", "skörda|VERB": "4", "såga|VERB": "4", "sökmotor|NOUN": "4", "drastiskt|ADV": "4", "dyrbar|ADJ": "4", "haka|VERB": "4", "knacka|VERB": "4", "offentlighet|NOUN": "4", "sekretess|NOUN": "4", "utkomma|VERB": "4", "indelning|NOUN": "4", "utomordentligt|ADV": "4", "olympisk|ADJ": "4", "skryta|VERB": "4", "ankomma|VERB": "4", "index|NOUN": "4", "umgänge|NOUN": "4", "välsignad|ADJ": "4", "avsky|VERB": "4", "förmoda|VERB": "4", "lyx|NOUN": "4", "skåp|NOUN": "4", "svamp|NOUN": "4", "uppehåll|NOUN": "4", "inbördes|ADJ": "4", "indikation|NOUN": "4", "jämlik|ADJ": "4", "staty|NOUN": "4", "uppförande|NOUN": "4", "överensstämmelse|NOUN": "4", "i grund och botten|ADV": "4", "puss|NOUN": "4", "spricka|NOUN": "4", "kemikalier|NOUN": "4", "konkurrenskraftig|ADJ": "4", "tankegång|NOUN": "4", "supporter|NOUN": "4", "symbolisk|ADJ": "4", "mervärde|NOUN": "4", "midsommar|NOUN": "4", "misstro|NOUN": "4", "fälla|NOUN": "4", "blues|NOUN": "4", "jury|NOUN": "4", "kör|NOUN": "4", "lyckligtvis|ADV": "4", "jordisk|ADJ": "4", "pumpa|VERB": "4", "harmoni|NOUN": "4", "trea|NOUN": "4", "avvägning|NOUN": "4", "markant|ADV": "4", "slopa|VERB": "4", "stål|NOUN": "4", "vinning|NOUN": "4", "främlingsfientlig|ADJ": "4", "mössa|NOUN": "4", "riksdagsman|NOUN": "4", "runtom|ADV": "4", "skikt|NOUN": "4", "avsevärd|ADJ": "4", "avvakta|VERB": "4", "dimma|NOUN": "4", "förundersökning|NOUN": "4", "huvudvärk|NOUN": "4", "ohälsa|NOUN": "4", "praktisera|VERB": "4", "rusta|VERB": "4", "subvention|NOUN": "4", "prisa|VERB": "4", "odemokratisk|ADJ": "4", "trilla|VERB": "4", "valfri|ADJ": "4", "mina|NOUN": "4", "ände|NOUN": "4", "hyresrätt|NOUN": "4", "härom|ADV": "4", "låga|NOUN": "4", "vital|ADJ": "4", "damm|NOUN": "4", "giftig|ADJ": "4", "pizza|NOUN": "4", "shopping|NOUN": "4", "färga|VERB": "4", "brygga|NOUN": "4", "kyckling|NOUN": "4", "löv|NOUN": "4", "specialist|NOUN": "4", "handlägga|VERB": "4", "hyckleri|NOUN": "4", "kännetecken|NOUN": "4", "överklass|NOUN": "4", "drivande|ADJ": "4", "arbetssätt|NOUN": "4", "hora|NOUN": "4", "nobelpris|NOUN": "4", "enkelhet|NOUN": "4", "förpliktelse|NOUN": "4", "larm|NOUN": "4", "lättnad|NOUN": "4", "predikan|NOUN": "4", "ammunition|NOUN": "4", "begär|NOUN": "4", "entydig|ADJ": "4", "missförstå|VERB": "4", "översvämning|NOUN": "4", "matcha|VERB": "4", "korrigera|VERB": "4", "försätta|VERB": "4", "frånvarande|ADJ": "4", "inblick|NOUN": "4", "ved|NOUN": "4", "mjukvara|NOUN": "4", "motpart|NOUN": "4", "riksdagsparti|NOUN": "4", "storskalig|ADJ": "4", "överflöd|NOUN": "4", "gröda|NOUN": "4", "jacka|NOUN": "4", "mottagande|NOUN": "4", "spårvagn|NOUN": "4", "återhämta|VERB": "4", "donera|VERB": "4", "sjukpenning|NOUN": "4", "bevarande|NOUN": "4", "bokhylla|NOUN": "4", "insida|NOUN": "4", "överraska|VERB": "4", "blöt|ADJ": "4", "relatera|VERB": "4", "underrättelsetjänst|NOUN": "4", "dynamik|NOUN": "4", "anmälning|NOUN": "4", "farhåga|NOUN": "4", "rovdjur|NOUN": "4", "tillsynsmyndighet|NOUN": "4", "adoptera|VERB": "4", "administrera|VERB": "4", "alltihop (vardagl. alltihopa)|PRON": "4", "dramatiskt|ADV": "4", "korkad|ADJ": "4", "marsch|NOUN": "4", "smäll|NOUN": "4", "less|ADJ": "4", "följande|ADJ": "4", "expedition|NOUN": "4", "heltäckande|ADJ": "4", "konvertera|VERB": "4", "i behov av|ADP": "4", "katastrofal|ADJ": "4", "näringsidkare|NOUN": "4", "otur|NOUN": "4", "flygning|NOUN": "4", "hierarki|NOUN": "4", "magasin|NOUN": "4", "plast|NOUN": "4", "stadig|ADJ": "4", "krävande|ADJ": "4", "täckt|ADJ": "4", "verifiera|VERB": "4", "blek|ADJ": "4", "förbjuden|ADJ": "4", "förnybar|ADJ": "4", "kyrkogård|NOUN": "4", "ovilja|NOUN": "4", "anarkist|NOUN": "4", "kartläggning|NOUN": "4", "krympa|VERB": "4", "skål|NOUN": "4", "underskatta|VERB": "4", "skifta|VERB": "4", "spänn|NOUN": "4", "auktion|NOUN": "4", "halka|VERB": "4", "kista|NOUN": "4", "sex|NOUN": "4", "vätska|NOUN": "4", "fascistisk|ADJ": "4", "hiss|NOUN": "4", "tå|NOUN": "4", "bestraffning|NOUN": "4", "bokstavligen|ADV": "4", "empirisk|ADJ": "4", "felaktigt|ADV": "4", "konfrontera|VERB": "4", "materia|NOUN": "4", "medborgerlig|ADJ": "4", "övergiven|ADJ": "4", "tillfredsställa|VERB": "4", "anmärkning|NOUN": "4", "nej|NOUN": "4", "skida|NOUN": "4", "förgäves|ADV": "4", "hiv|NOUN": "4", "kabel|NOUN": "4", "projektledare|NOUN": "4", "strikt|ADV": "4", "klinik|NOUN": "4", "råtta|NOUN": "4", "strömning|NOUN": "4", "kandidera|VERB": "4", "revolutionär|NOUN": "4", "ritning|NOUN": "4", "utmed|ADP": "4", "visdom|NOUN": "4", "uppfostra|VERB": "4", "lagändring|NOUN": "4", "så länge (som)|SCONJ": "4", "kulturarv|NOUN": "4", "nordlig|ADJ": "4", "plantera|VERB": "4", "chaufför|NOUN": "4", "inuti|ADP": "4", "förbruka|VERB": "4", "budgetproposition|NOUN": "4", "ceremoni|NOUN": "4", "uran|NOUN": "4", "aktualisera|VERB": "4", "barnfamilj|NOUN": "4", "population|NOUN": "4", "undanröja|VERB": "4", "utväg|NOUN": "4", "entreprenörskap|NOUN": "4", "godtagbar|ADJ": "4", "mardröm|NOUN": "4", "storebror|NOUN": "4", "isolera|VERB": "4", "kalas|NOUN": "4", "kopiering|NOUN": "4", "paroll|NOUN": "4", "shoppa|VERB": "4", "språkbruk|NOUN": "4", "diabetes|NOUN": "4", "fortlöpande|ADJ": "4", "klädsel|NOUN": "4", "svagt|ADV": "4", "ämbete|NOUN": "4", "historik|NOUN": "4", "intyg|NOUN": "4", "konversation|NOUN": "4", "växel|NOUN": "4", "byråkratisk|ADJ": "4", "etablering|NOUN": "4", "förnuftig|ADJ": "4", "hedra|VERB": "4", "omedveten|ADJ": "4", "stundtals|ADV": "4", "tjata|VERB": "4", "tjeckisk|ADJ": "4", "åtanke|NOUN": "4", "fördelaktig|ADJ": "4", "assistent|NOUN": "4", "läskig|ADJ": "4", "nationalekonomi|NOUN": "4", "återfå|VERB": "4", "övernaturlig|ADJ": "4", "elektricitet|NOUN": "4", "grovt|ADV": "4", "javisst (el. ja visst)|INTJ": "4", "beskylla|VERB": "4", "obegränsad|ADJ": "4", "anordning|NOUN": "4", "fluga|NOUN": "4", "förråd|NOUN": "4", "spänna|VERB": "4", "oönskad|ADJ": "4", "marschera|VERB": "4", "päls|NOUN": "4", "till vara|ADV": "4", "slant|NOUN": "4", "upprättande|NOUN": "4", "överdriva|VERB": "4", "reparera|VERB": "4", "central|NOUN": "4", "erövring|NOUN": "4", "justering|NOUN": "4", "nedanstående|ADJ": "4", "propagera|VERB": "4", "talesman|NOUN": "4", "uppträdande|NOUN": "4", "tandläkare|NOUN": "4", "utförande|NOUN": "4", "utgivare|NOUN": "4", "underordnad|ADJ": "4", "explosion|NOUN": "4", "fraktion|NOUN": "4", "renovera|VERB": "4", "snyggt|ADV": "4", "beröva|VERB": "4", "japan|NOUN": "4", "omvandling|NOUN": "4", "tillåtelse|NOUN": "4", "vidrig|ADJ": "4", "förmögen|ADJ": "4", "nedanför|ADP": "4", "oförmögen|ADJ": "4", "slösa|VERB": "4", "arbetsmarknadspolitik|NOUN": "4", "inkomstskatt|NOUN": "4", "skämta|VERB": "4", "underrätta|VERB": "4", "världslig|ADJ": "4", "cigarett|NOUN": "4", "hälsosam|ADJ": "4", "skalle|NOUN": "4", "spädbarn|NOUN": "4", "domslut|NOUN": "4", "dyrka|VERB": "4", "utmärkelse|NOUN": "4", "katalog|NOUN": "4", "bredband|NOUN": "4", "kemi|NOUN": "4", "foster|NOUN": "5", "tillfällighet|NOUN": "5", "enastående|ADJ": "5", "rökning|NOUN": "5", "trots|NOUN": "5", "muta|NOUN": "5", "motgång|NOUN": "5", "människosyn|NOUN": "5", "omvända|VERB": "5", "sammanbrott|NOUN": "5", "auktoritär|ADJ": "5", "bebis|NOUN": "5", "fat|NOUN": "5", "hunger|NOUN": "5", "metafor|NOUN": "5", "understödja|VERB": "5", "anamma|VERB": "5", "arrestera|VERB": "5", "barriär|NOUN": "5", "best|NOUN": "5", "fästning|NOUN": "5", "immateriell|ADJ": "5", "vansinne|NOUN": "5", "involvera|VERB": "5", "hopplös|ADJ": "5", "införliva|VERB": "5", "tacksamhet|NOUN": "5", "återkalla|VERB": "5", "jämnt|ADJ": "5", "extremist|NOUN": "5", "civilbefolkning|NOUN": "5", "förtvivlan|NOUN": "5", "löntagare|NOUN": "5", "åratal|NOUN": "5", "överträffa|VERB": "5", "flitig|ADJ": "5", "härleda|VERB": "5", "greve|NOUN": "5", "internt|ADV": "5", "soppa|NOUN": "5", "tvivelaktig|ADJ": "5", "ändamålsenlig|ADJ": "5", "byråkrat|NOUN": "5", "lagstiftande|ADJ": "5", "civiliserad|ADJ": "5", "fjäll|NOUN": "5", "knäcka|VERB": "5", "likgiltig|ADJ": "5", "nationalist|NOUN": "5", "offensiv|ADJ": "5", "socialbidrag|NOUN": "5", "befästa|VERB": "5", "väninna|NOUN": "5", "blixt|NOUN": "5", "bevisligen|ADV": "5", "fräsch|ADJ": "5", "ivrig|ADJ": "5", "mus|NOUN": "5", "tillkännagivande|NOUN": "5", "lojal|ADJ": "5", "småföretag|NOUN": "5", "terapi|NOUN": "5", "undanta|VERB": "5", "frekvens|NOUN": "5", "givande|ADJ": "5", "i ljuset av|ADP": "5", "komisk|ADJ": "5", "kostnadsfri|ADJ": "5", "uniform|NOUN": "5", "utfrågning|NOUN": "5", "godhet|NOUN": "5", "tysta|VERB": "5", "bombning|NOUN": "5", "engelskspråkig|ADJ": "5", "beslag|NOUN": "5", "vapenvila|NOUN": "5", "buller|NOUN": "5", "intervention|NOUN": "5", "lagring|NOUN": "5", "utbyta|VERB": "5", "svin|NOUN": "5", "lagom|ADJ": "5", "doktrin|NOUN": "5", "klick|NOUN": "5", "stämpla|VERB": "5", "uppfostran|NOUN": "5", "bilateral|ADJ": "5", "bostadsrätt|NOUN": "5", "iakttagelse|NOUN": "5", "på sistone|ADV": "5", "påskynda|VERB": "5", "sponsra|VERB": "5", "avbrott|NOUN": "5", "bestånd|NOUN": "5", "hantverkare|NOUN": "5", "sjukskrivning|NOUN": "5", "slakta|VERB": "5", "uppröra|VERB": "5", "besittning|NOUN": "5", "fasa|NOUN": "5", "konfrontation|NOUN": "5", "trådlös|ADJ": "5", "pub|NOUN": "5", "biverkning|NOUN": "5", "dragning|NOUN": "5", "logiskt|ADV": "5", "österut|ADV": "5", "deckare|NOUN": "5", "dåtid|NOUN": "5", "cynisk|ADJ": "5", "poetisk|ADJ": "5", "kostsam|ADJ": "5", "misslyckad|ADJ": "5", "prioritet|NOUN": "5", "fascist|NOUN": "5", "frestelse|NOUN": "5", "trösta|VERB": "5", "uppriktigt|ADV": "5", "världsekonomi|NOUN": "5", "summera|VERB": "5", "fängelsestraff|NOUN": "5", "invigning|NOUN": "5", "revisor|NOUN": "5", "samisk|ADJ": "5", "så snart som|ADV": "5", "underminera|VERB": "5", "medgivande|NOUN": "5", "tvätt|NOUN": "5", "guvernör|NOUN": "5", "adekvat|ADJ": "5", "brottas|VERB": "5", "hantverk|NOUN": "5", "minus|ADV": "5", "fullborda|VERB": "5", "latinsk|ADJ": "5", "stabilisera|VERB": "5", "kvantitet|NOUN": "5", "huvudroll|NOUN": "5", "hög|NOUN": "5", "knepig|ADJ": "5", "överblick|NOUN": "5", "berömma|VERB": "5", "räckvidd|NOUN": "5", "utifrån|ADV": "5", "västlig|ADJ": "5", "skicklighet|NOUN": "5", "bestraffa|VERB": "5", "spik|NOUN": "5", "akademiker|NOUN": "5", "författarskap|NOUN": "5", "närvara|VERB": "5", "sola|VERB": "5", "association|NOUN": "5", "exil|NOUN": "5", "förbehåll|NOUN": "5", "hämma|VERB": "5", "nominera|VERB": "5", "viska|VERB": "5", "koalition|NOUN": "5", "spektakulär|ADJ": "5", "teoretiskt|ADV": "5", "handfull|NOUN": "5", "ugn|NOUN": "5", "geografi|NOUN": "5", "meditation|NOUN": "5", "betoning|NOUN": "5", "brevlåda|NOUN": "5", "förfoga|VERB": "5", "heja|VERB": "5", "ironisk|ADJ": "5", "skrivare|NOUN": "5", "valdeltagande|NOUN": "5", "lamm|NOUN": "5", "berika|VERB": "5", "brytning|NOUN": "5", "flyktingpolitik|NOUN": "5", "porr|NOUN": "5", "flöda|VERB": "5", "revolt|NOUN": "5", "snällt|ADV": "5", "vika|ADV": "5", "ekosystem|NOUN": "5", "heterosexuell|ADJ": "5", "kolumn|NOUN": "5", "lyssnare|NOUN": "5", "möjligt|ADV": "5", "utebli|VERB": "5", "underkasta|VERB": "5", "salong|NOUN": "5", "sjöfart|NOUN": "5", "tapet|NOUN": "5", "bråttom|ADV": "5", "kraftverk|NOUN": "5", "spotta|VERB": "5", "duscha|VERB": "5", "attrahera|VERB": "5", "måste|NOUN": "5", "ovannämnd|ADJ": "5", "tänkare|NOUN": "5", "morot|NOUN": "5", "censurera|VERB": "5", "lagtext|NOUN": "5", "lindra|VERB": "5", "vilse|ADV": "5", "förenkling|NOUN": "5", "tolerera|VERB": "5", "löst|ADV": "5", "sankt (förk. s:t)|ADJ": "5", "överflödig|ADJ": "5", "omnämna|VERB": "5", "pund|NOUN": "5", "slöseri|NOUN": "5", "formel|NOUN": "5", "drink|NOUN": "5", "förväntan|NOUN": "5", "lunga|NOUN": "5", "vårdcentral|NOUN": "5", "ödmjukhet|NOUN": "5", "överdrift|NOUN": "5", "häpnadsväckande|ADJ": "5", "urskilja|VERB": "5", "frigörelse|NOUN": "5", "monetär|ADJ": "5", "tobak|NOUN": "5", "tråkigt|ADV": "5", "förordna|VERB": "5", "femma|NOUN": "5", "livslängd|NOUN": "5", "sval|ADJ": "5", "telefonnummer|NOUN": "5", "analytiker|NOUN": "5", "avspegla|VERB": "5", "psykiatrisk|ADJ": "5", "rebell|NOUN": "5", "droppa|VERB": "5", "tugga|VERB": "5", "kval|NOUN": "5", "läroplan|NOUN": "5", "psalm|NOUN": "5", "sårbar|ADJ": "5", "kår|NOUN": "5", "luthersk|ADJ": "5", "stel|ADJ": "5", "tydliggöra|VERB": "5", "barnslig|ADJ": "5", "betraktelse|NOUN": "5", "fortgå|VERB": "5", "optimistisk|ADJ": "5", "tillfredsställelse|NOUN": "5", "välmående|ADJ": "5", "applicera|VERB": "5", "förkortning|NOUN": "5", "jämställa|VERB": "5", "runt omkring|ADV": "5", "välsigna|VERB": "5", "donation|NOUN": "5", "laddad|ADJ": "5", "monument|NOUN": "5", "blomma|VERB": "5", "hona|NOUN": "5", "prick|NOUN": "5", "humanistisk|ADJ": "5", "intressent|NOUN": "5", "parameter|NOUN": "5", "sopa|VERB": "5", "streck|NOUN": "5", "ikon|NOUN": "5", "insekt|NOUN": "5", "dotterbolag|NOUN": "5", "irakier|NOUN": "5", "istid|NOUN": "5", "till slut|ADV": "5", "försening|NOUN": "5", "färja|NOUN": "5", "förståelig|ADJ": "5", "prenumerera|VERB": "5", "ansluten|ADJ": "5", "romantik|NOUN": "5", "bisarr|ADJ": "5", "förfalla|VERB": "5", "lås|NOUN": "5", "principiellt|ADV": "5", "samförstånd|NOUN": "5", "jazz|NOUN": "5", "ritual|NOUN": "5", "segel|NOUN": "5", "exotisk|ADJ": "5", "informationssamhälle|NOUN": "5", "lukt|NOUN": "5", "skrapa|VERB": "5", "uppgradera|VERB": "5", "mäklare|NOUN": "5", "reservera|VERB": "5", "bur|NOUN": "5", "snöa|VERB": "5", "anteckna|VERB": "5", "box|NOUN": "5", "korsning|NOUN": "5", "legitimera|VERB": "5", "förfärlig|ADJ": "5", "förvånansvärt|ADV": "5", "kretsa|VERB": "5", "implementera|VERB": "5", "alster|NOUN": "5", "energikälla|NOUN": "5", "livsfarlig|ADJ": "5", "livskvalitet|NOUN": "5", "måttlig|ADJ": "5", "tryggt|ADV": "5", "bäck|NOUN": "5", "förtal|NOUN": "5", "förutsägbar|ADJ": "5", "intensifiera|VERB": "5", "naturresurs|NOUN": "5", "otänkbar|ADJ": "5", "varsel|NOUN": "5", "tillbehör|NOUN": "5", "betong|NOUN": "5", "nybörjare|NOUN": "5", "ruin|NOUN": "5", "sortiment|NOUN": "5", "nyans|NOUN": "5", "uppbära|VERB": "5", "arkeologisk|ADJ": "5", "okunnighet|NOUN": "5", "anseende|NOUN": "5", "förbannelse|NOUN": "5", "jubla|VERB": "5", "lejon|NOUN": "5", "session|NOUN": "5", "effektivisera|VERB": "5", "hotfull|ADJ": "5", "miljöpolitik|NOUN": "5", "storföretag|NOUN": "5", "suveränitet|NOUN": "5", "utanför|ADV": "5", "landshövding|NOUN": "5", "statsbidrag|NOUN": "5", "storslagen|ADJ": "5", "separera|VERB": "5", "firande|NOUN": "5", "hyllning|NOUN": "5", "oljepris|NOUN": "5", "biologi|NOUN": "5", "rimligtvis|ADV": "5", "arbetarparti|NOUN": "5", "beskåda|VERB": "5", "briljant|ADJ": "5", "lott|NOUN": "5", "kidnappa|VERB": "5", "girighet|NOUN": "5", "härröra|VERB": "5", "på sätt och vis|ADV": "5", "framlägga|VERB": "5", "förorsaka|VERB": "5", "häck|NOUN": "5", "hemvist|NOUN": "5", "andetag|NOUN": "5", "berusad|ADJ": "5", "tortera|VERB": "5", "kanadensisk|ADJ": "5", "protestantisk|ADJ": "5", "läktare|NOUN": "5", "marxist|NOUN": "5", "peta|VERB": "5", "sakkunnig|ADJ": "5", "svängning|NOUN": "5", "tanka|VERB": "5", "sympatisk|ADJ": "5", "översikt|NOUN": "5", "midnatt|NOUN": "5", "amatör|NOUN": "5", "befalla|VERB": "5", "handledare|NOUN": "5", "bostadsmarknad|NOUN": "5", "klappa|VERB": "5", "media|NOUN": "5", "när som helst|ADV": "5", "pil|NOUN": "5", "rättsstat|NOUN": "5", "röra|NOUN": "5", "vålla|VERB": "5", "blygsam|ADJ": "5", "exponering|NOUN": "5", "närområde|NOUN": "5", "otrogen|ADJ": "5", "varva|VERB": "5", "regent|NOUN": "5", "bunt|NOUN": "5", "fostra|VERB": "5", "funktionell|ADJ": "5", "klinisk|ADJ": "5", "värdegrund|NOUN": "5", "förutsäga|VERB": "5", "begrunda|VERB": "5", "tennis|NOUN": "5", "destination|NOUN": "5", "taktisk|ADJ": "5", "österrikisk|ADJ": "5", "manifestera|VERB": "5", "förakta|VERB": "5", "invandringspolitik|NOUN": "5", "utbrista|VERB": "5", "aids|NOUN": "5", "bekanta|VERB": "5", "utövare|NOUN": "5", "angå|VERB": "5", "förlossning|NOUN": "5", "återgång|NOUN": "5", "procedur|NOUN": "5", "äventyra|VERB": "5", "rep|NOUN": "5", "sväva|VERB": "5", "diet|NOUN": "5", "filter|NOUN": "5", "gratis|ADJ": "5", "legendarisk|ADJ": "5", "plagg|NOUN": "5", "impuls|NOUN": "5", "parkering|NOUN": "5", "beståndsdel|NOUN": "5", "brottslig|ADJ": "5", "årstid|NOUN": "5", "underlåta|VERB": "5", "episod|NOUN": "5", "kock|NOUN": "5", "affärsman|NOUN": "5", "högkonjunktur|NOUN": "5", "lur|NOUN": "5", "nu|NOUN": "5", "opinionsbildning|NOUN": "5", "premiss|NOUN": "5", "insistera|VERB": "5", "grafik|NOUN": "5", "munk|NOUN": "5", "skörd|NOUN": "5", "dräkt|NOUN": "5", "galenskap|NOUN": "5", "franska|NOUN": "5", "pistol|NOUN": "5", "pyssla|VERB": "5", "urholka|VERB": "5", "galning|NOUN": "5", "hugg|NOUN": "5", "preferens|NOUN": "5", "uppslag|NOUN": "5", "exploatera|VERB": "5", "förväxla|VERB": "5", "tomat|NOUN": "5", "ocean|NOUN": "5", "cyklist|NOUN": "5", "näve|NOUN": "5", "omstrukturering|NOUN": "5", "restriktiv|ADJ": "5", "skina|VERB": "5", "skulptur|NOUN": "5", "ättling|NOUN": "5", "helgon|NOUN": "5", "utstå|VERB": "5", "envisas|VERB": "5", "pedagogik|NOUN": "5", "postning|NOUN": "5", "trygga|VERB": "5", "uppmärksam|ADJ": "5", "bädda|VERB": "5", "fuktig|ADJ": "5", "fundament|NOUN": "5", "reformation|NOUN": "5", "grilla|VERB": "5", "italienare|NOUN": "5", "famn|NOUN": "5", "genomgripande|ADJ": "5", "skägg|NOUN": "5", "slappna|VERB": "5", "medalj|NOUN": "5", "expansiv|ADJ": "5", "matlagning|NOUN": "5", "rytm|NOUN": "5", "elefant|NOUN": "5", "patetisk|ADJ": "5", "batteri|NOUN": "5", "tippa|VERB": "5", "ambulans|NOUN": "5", "bearbetning|NOUN": "5", "huvudkontor|NOUN": "5", "precisera|VERB": "5", "folkmassa|NOUN": "5", "ohållbar|ADJ": "5", "revision|NOUN": "5", "såra|VERB": "5", "mix|NOUN": "5", "vy|NOUN": "5", "diplomat|NOUN": "5", "affisch|NOUN": "5", "associera|VERB": "5", "kalkyl|NOUN": "5", "konstgjord|ADJ": "5", "polack|NOUN": "5", "renovering|NOUN": "5", "maffia|NOUN": "5", "snickare|NOUN": "5", "teolog|NOUN": "5", "väster om|ADP": "5", "kontinuitet|NOUN": "5", "marginell|ADJ": "5", "ojämn|ADJ": "5", "skoja|VERB": "5", "tangentbord|NOUN": "5", "migration|NOUN": "5", "säck|NOUN": "5", "körning|NOUN": "5", "blond|ADJ": "5", "dygd|NOUN": "5", "förorening|NOUN": "5", "svenskspråkig|ADJ": "5", "lera|NOUN": "5", "befattning|NOUN": "5", "föredöme|NOUN": "5", "genetiskt|ADV": "5", "sucka|VERB": "5", "framhäva|VERB": "5", "laboratorium|NOUN": "5", "strypa|VERB": "5", "kroppslig|ADJ": "5", "pool|NOUN": "5", "sionism|NOUN": "5", "uttag|NOUN": "5", "begynnelse|NOUN": "5", "likartad|ADJ": "5", "slakt|NOUN": "5", "naturvetenskap|NOUN": "5", "premie|NOUN": "5", "snus|NOUN": "5", "tillgå|VERB": "5", "vadå|INTJ": "5", "valresultat|NOUN": "5", "västerut|ADV": "5", "diamant|NOUN": "5", "kulle|NOUN": "5", "avlyssna|VERB": "5", "bärbar|ADJ": "5", "förkylning|NOUN": "5", "piano|NOUN": "5", "plåga|NOUN": "5", "signalera|VERB": "5", "snubbe|NOUN": "5", "eftergift|NOUN": "5", "major|NOUN": "5", "veterinär|NOUN": "5", "utopi|NOUN": "5", "författa|VERB": "5", "gräsmatta|NOUN": "5", "bifoga|VERB": "5", "parkera|VERB": "5", "fastland|NOUN": "5", "mentalitet|NOUN": "5", "slagfält|NOUN": "5", "stimulans|NOUN": "5", "proffs|NOUN": "5", "ekvation|NOUN": "5", "repris|NOUN": "5", "rådgivande|ADJ": "5", "vinnande|ADJ": "5", "diskret|ADJ": "5", "befallning|NOUN": "5", "pipa|NOUN": "5", "kjol|NOUN": "5", "bubbla|NOUN": "5", "mirakel|NOUN": "5", "hednisk|ADJ": "5", "lök|NOUN": "5", "infektion|NOUN": "5", "integrering|NOUN": "5", "uträtta|VERB": "5", "älskling|NOUN": "5", "pedagog|NOUN": "5", "kvalitativ|ADJ": "5", "motorcykel|NOUN": "5", "styrelseledamot|NOUN": "5", "tvärt|ADV": "5", "domän|NOUN": "5", "subjekt|NOUN": "5", "fana|NOUN": "5", "fax|NOUN": "6", "belasta|VERB": "5", "föreläsare|NOUN": "5", "lagstiftare|NOUN": "5", "högkvarter|NOUN": "5", "fascinera|VERB": "5", "fånig|ADJ": "5", "administratör|NOUN": "5", "förälskad|ADJ": "5", "gagna|VERB": "5", "modifiera|VERB": "5", "realisera|VERB": "5", "samlag|NOUN": "5", "skymta|VERB": "5", "utbredning|NOUN": "5", "utkant|NOUN": "5", "envis|ADJ": "5", "syndare|NOUN": "5", "paradox|NOUN": "5", "bräda|NOUN": "5", "ordbok|NOUN": "5", "översättare|NOUN": "5", "avkomma|NOUN": "5", "avlägga|VERB": "5", "utnämning|NOUN": "5", "riddare|NOUN": "5", "handikapp|NOUN": "5", "myra|NOUN": "5", "hop|NOUN": "5", "föreläsa|VERB": "5", "besläktad|ADJ": "5", "halvö|NOUN": "5", "sammanslagning|NOUN": "5", "yngling|NOUN": "5", "klassificera|VERB": "5", "spruta|VERB": "5", "spärra|VERB": "5", "biograf|NOUN": "5", "klan|NOUN": "5", "löpning|NOUN": "5", "profit|NOUN": "5", "hållbarhet|NOUN": "5", "foder|NOUN": "5", "framsida|NOUN": "5", "solidarisk|ADJ": "5", "tallrik|NOUN": "5", "nominering|NOUN": "5", "handbok|NOUN": "5", "debut|NOUN": "5", "försiktighet|NOUN": "5", "groda|NOUN": "5", "hobby|NOUN": "5", "bidragande|ADJ": "5", "blomstra|VERB": "5", "välbefinnande|NOUN": "5", "deg|NOUN": "5", "demo|NOUN": "5", "fiskare|NOUN": "5", "ryggsäck|NOUN": "5", "behaga|VERB": "5", "ekumenisk|ADJ": "5", "partikel|NOUN": "5", "svettig|ADJ": "5", "tårta|NOUN": "5", "utsida|NOUN": "5", "drunkna|VERB": "5", "kognitiv|ADJ": "5", "prägel|NOUN": "5", "klang|NOUN": "5", "pc|NOUN": "5", "faktura|NOUN": "5", "oroväckande|ADJ": "5", "broschyr|NOUN": "5", "mästerskap|NOUN": "5", "terror|NOUN": "5", "duk|NOUN": "5", "expertis|NOUN": "5", "jungfru|NOUN": "5", "utgivning|NOUN": "5", "avundsjuka|NOUN": "5", "multinationell|ADJ": "5", "vett|NOUN": "5", "insättning|NOUN": "5", "statisk|ADJ": "5", "stavning|NOUN": "5", "steka|VERB": "5", "bedra|VERB": "5", "förvandling|NOUN": "5", "snäv|ADJ": "5", "läka|VERB": "5", "nagel|NOUN": "5", "utdragen|ADJ": "5", "överordnad|ADJ": "5", "tillbe|VERB": "5", "avsändare|NOUN": "5", "beklaglig|ADJ": "5", "sköld|NOUN": "5", "syre|NOUN": "5", "bubbla|VERB": "5", "kväva|VERB": "5", "motstå|VERB": "5", "väktare|NOUN": "5", "express|NOUN": "5", "häxa|NOUN": "5", "irritera|VERB": "5", "lärobok|NOUN": "5", "nerv|NOUN": "5", "pendla|VERB": "5", "trakassera|VERB": "5", "förvaring|NOUN": "5", "oskuld|NOUN": "5", "sydlig|ADJ": "5", "gudinna|NOUN": "5", "sponsor|NOUN": "5", "bekantskap|NOUN": "5", "skoj|ADJ": "5", "filial|NOUN": "5", "kvalifikation|NOUN": "5", "ratificera|VERB": "5", "spis|NOUN": "5", "strumpa|NOUN": "5", "hetta|NOUN": "5", "kyssa|VERB": "5", "sekundär|ADJ": "5", "utmanande|ADJ": "5", "avbilda|VERB": "5", "segling|NOUN": "5", "drastisk|ADJ": "5", "korg|NOUN": "5", "avsiktligt|ADV": "5", "tystna|VERB": "5", "underjordisk|ADJ": "5", "entusiastisk|ADJ": "5", "talarstol|NOUN": "5", "omöjlighet|NOUN": "5", "kriga|VERB": "5", "kylskåp|NOUN": "5", "skoj|NOUN": "5", "omkomma|VERB": "5", "territoriell|ADJ": "5", "provisorisk|ADJ": "5", "tablett|NOUN": "5", "galax|NOUN": "5", "sallad|NOUN": "5", "berömd|ADJ": "5", "hjälm|NOUN": "5", "teknologisk|ADJ": "5", "försumma|VERB": "5", "föråldrad|ADJ": "5", "komplexitet|NOUN": "5", "kronisk|ADJ": "5", "geni|NOUN": "5", "kvadratmeter|NOUN": "5", "tillfoga|VERB": "5", "upprepning|NOUN": "5", "cirkulera|VERB": "5", "kvantitativ|ADJ": "5", "kvot|NOUN": "5", "hallå|INTJ": "5", "tröskel|NOUN": "5", "syndrom|NOUN": "5", "tvilling|NOUN": "5", "modernisera|VERB": "5", "stämpel|NOUN": "5", "autonomi|NOUN": "5", "mjöl|NOUN": "5", "vägledande|ADJ": "5", "slagsmål|NOUN": "5", "semifinal|NOUN": "5", "diktera|VERB": "5", "lärorik|ADJ": "5", "samarbetspartner|NOUN": "5", "envar|PRON": "5", "bokhandel|NOUN": "5", "dunkel|ADJ": "5", "reparation|NOUN": "5", "docka|NOUN": "5", "obehag|NOUN": "5", "originell|ADJ": "5", "galleri|NOUN": "5", "ökänd|ADJ": "5", "mottagning|NOUN": "5", "intensitet|NOUN": "5", "modernisering|NOUN": "5", "visuell|ADJ": "5", "kommentator|NOUN": "5", "beskydd|NOUN": "5", "döv|ADJ": "5", "knäppa|VERB": "5", "grundlig|ADJ": "5", "husdjur|NOUN": "5", "halvvägs|ADV": "5", "tomhet|NOUN": "5", "ansats|NOUN": "5", "iskall|ADJ": "5", "ofattbar|ADJ": "5", "tiger|NOUN": "5", "applikation|NOUN": "5", "självstyre|NOUN": "5", "mästerverk|NOUN": "5", "svett|NOUN": "5", "studsa|VERB": "5", "optimism|NOUN": "5", "uppgradering|NOUN": "5", "befordra|VERB": "5", "intyga|VERB": "5", "vinka|VERB": "5", "motsägelse|NOUN": "5", "martyr|NOUN": "5", "satellit|NOUN": "5", "uppriktig|ADJ": "5", "bedrift|NOUN": "5", "förvaltare|NOUN": "5", "biträdande|ADJ": "5", "segrare|NOUN": "5", "dumpa|VERB": "5", "övervikt|NOUN": "5", "kollapsa|VERB": "5", "städning|NOUN": "5", "borra|VERB": "5", "nyfödd|ADJ": "5", "smink|NOUN": "5", "parentes|NOUN": "5", "infödd|ADJ": "5", "irritation|NOUN": "5", "rutten|ADJ": "5", "fakultet|NOUN": "5", "skiss|NOUN": "5", "rand|NOUN": "5", "festa|VERB": "5", "frekvent|ADJ": "5", "prestanda|NOUN": "5", "djärv|ADJ": "5", "omtyckt|ADJ": "5", "skrik|NOUN": "5", "förtvivlad|ADJ": "5", "uttrycklig|ADJ": "5", "signera|VERB": "5", "experimentera|VERB": "5", "födsel|NOUN": "5", "ombyggnad|NOUN": "5", "avgrund|NOUN": "5", "kapell|NOUN": "5", "planta|NOUN": "5", "våt|ADJ": "5", "fångenskap|NOUN": "5", "korrekthet|NOUN": "5", "variabel|NOUN": "5", "formulär|NOUN": "5", "gap|NOUN": "5", "manifest|NOUN": "5", "handlare|NOUN": "5", "mobilisering|NOUN": "5", "återförsäljare|NOUN": "5", "fördjupning|NOUN": "5", "räv|NOUN": "5", "anvisa|VERB": "5", "definitiv|ADJ": "5", "misstänksam|ADJ": "5", "intervall|NOUN": "5", "gryta|NOUN": "5", "återvinna|VERB": "5", "frakta|VERB": "5", "gumma|NOUN": "5", "ojämlikhet|NOUN": "5", "krut|NOUN": "5", "precision|NOUN": "5", "anslå|VERB": "5", "orealistisk|ADJ": "5", "copyright|NOUN": "5", "företräde|NOUN": "5", "minimum|NOUN": "5", "skolgång|NOUN": "5", "giltighet|NOUN": "5", "anknyta|VERB": "5", "avskeda|VERB": "5", "barmhärtighet|NOUN": "5", "gevär|NOUN": "5", "visum|NOUN": "5", "analytisk|ADJ": "5", "intrig|NOUN": "5", "förkorta|VERB": "5", "påträffa|VERB": "5", "skådespel|NOUN": "5", "avtryck|NOUN": "5", "disponera|VERB": "5", "knuffa|VERB": "5", "vägran|NOUN": "5", "charm|NOUN": "5", "uthärda|VERB": "5", "högtidlig|ADJ": "5", "komplikation|NOUN": "5", "delegat|NOUN": "5", "socialförsäkring|NOUN": "5", "öm|ADJ": "5", "bälte|NOUN": "5", "privatisera|VERB": "5", "lillebror|NOUN": "5", "smuts|NOUN": "5", "kudde|NOUN": "5", "slätt|NOUN": "5", "kondom|NOUN": "5", "tank|NOUN": "5", "bråkdel|NOUN": "5", "ögonbryn|NOUN": "5", "undkomma|VERB": "5", "hejdå (el. hej då)|INTJ": "5", "spannmål|NOUN": "5", "uttal|NOUN": "5", "kompositör|NOUN": "5", "korn|NOUN": "5", "täckning|NOUN": "5", "anstalt|NOUN": "5", "förmedling|NOUN": "5", "deprimerad|ADJ": "5", "sammankomst|NOUN": "5", "vänligen|ADV": "5", "grymhet|NOUN": "5", "nykter|ADJ": "5", "solid|ADJ": "5", "idealisk|ADJ": "5", "pyramid|NOUN": "5", "stövel|NOUN": "5", "gråt|NOUN": "5", "täcke|NOUN": "5", "blinka|VERB": "5", "gränd|NOUN": "5", "otillåten|ADJ": "5", "prestige|NOUN": "5", "tolk|NOUN": "5", "reträtt|NOUN": "5", "nolla|NOUN": "5", "bricka|NOUN": "5", "korrigering|NOUN": "5", "lyxig|ADJ": "5", "reaktor|NOUN": "5", "banan|NOUN": "5", "kult|NOUN": "5", "komedi|NOUN": "5", "trick|NOUN": "5", "separation|NOUN": "5", "avlösa|VERB": "5", "betvivla|VERB": "5", "likaledes|ADV": "5", "retur|NOUN": "5", "dussin|NOUN": "5", "kylig|ADJ": "5", "dröjsmål|NOUN": "5", "grädde|NOUN": "5", "intellekt|NOUN": "5", "aggression|NOUN": "5", "buske|NOUN": "5", "minderårig|ADJ": "5", "spinna|VERB": "5", "interaktion|NOUN": "5", "terminologi|NOUN": "5", "östlig|ADJ": "5", "avsked|NOUN": "5", "hal|ADJ": "5", "rival|NOUN": "5", "proklamera|VERB": "5", "sofistikerad|ADJ": "5", "spruta|NOUN": "5", "anständig|ADJ": "5", "pump|NOUN": "5", "sexig|ADJ": "5", "förflyttning|NOUN": "5", "huvudsak|NOUN": "5", "utelämna|VERB": "5", "boskap|NOUN": "5", "exponera|VERB": "5", "lila|ADJ": "5", "tillägna|VERB": "5", "genus|NOUN": "5", "verb|NOUN": "5", "köpman|NOUN": "5", "vidarebefordra|VERB": "5", "frånta|VERB": "5", "interaktiv|ADJ": "5", "lagstifta|VERB": "5", "specialitet|NOUN": "5", "stråla|VERB": "5", "domkyrka|NOUN": "5", "slapp|ADJ": "5", "utvinna|VERB": "5", "upphöjd|ADJ": "5", "vykort|NOUN": "5", "assistans|NOUN": "5", "begåvning|NOUN": "5", "måleri|NOUN": "5", "påhitt|NOUN": "5", "kompakt|ADJ": "5", "samtycka|VERB": "5", "hälsovård|NOUN": "5", "lyft|NOUN": "5", "asfalt|NOUN": "5", "underkänna|VERB": "5", "uppoffring|NOUN": "5", "utrusta|VERB": "5", "förflyta|VERB": "5", "handledning|NOUN": "5", "oenighet|NOUN": "5", "slogan|NOUN": "5", "triumf|NOUN": "5", "färdigställa|VERB": "5", "skötsel|NOUN": "5", "portal|NOUN": "5", "överdrivet|ADV": "5", "applådera|VERB": "5", "husvagn|NOUN": "5", "vodka|NOUN": "5", "lansering|NOUN": "5", "handduk|NOUN": "5", "honung|NOUN": "5", "kanin|NOUN": "5", "målare|NOUN": "5", "plågsam|ADJ": "5", "trollkarl|NOUN": "5", "avancera|VERB": "5", "homogen|ADJ": "5", "skingra|VERB": "5", "underordna|VERB": "5", "överlägsenhet|NOUN": "5", "krocka|VERB": "5", "filt|NOUN": "5", "herravälde|NOUN": "5", "ryttare|NOUN": "5", "peppar|NOUN": "5", "nominell|ADJ": "5", "spola|VERB": "5", "defensiv|ADJ": "5", "katedral|NOUN": "5", "fjärran|ADJ": "5", "skär|ADJ": "5", "desperation|NOUN": "5", "blöda|VERB": "5", "ört|NOUN": "5", "avslappnad|ADJ": "5", "efterlevnad|NOUN": "5", "resande|NOUN": "5", "bär|NOUN": "5", "mysterium|NOUN": "5", "omvänt|ADV": "5", "lillasyster|NOUN": "5", "massage|NOUN": "5", "märkbar|ADJ": "5", "hane|NOUN": "5", "regelrätt|ADJ": "5", "gryning|NOUN": "5", "gudom|NOUN": "5", "överste|NOUN": "5", "uttråkad|ADJ": "5", "helikopter|NOUN": "5", "parasit|NOUN": "5", "utgrävning|NOUN": "5", "drake|NOUN": "5", "kryssa|VERB": "5", "stolpe|NOUN": "5", "kartong|NOUN": "5", "realism|NOUN": "5", "stackare|NOUN": "5", "höft|NOUN": "5", "skinka|NOUN": "5", "stökig|ADJ": "5", "råna|VERB": "5", "anförtro|VERB": "5", "försäljare|NOUN": "5", "gränssnitt|NOUN": "5", "stängning|NOUN": "5", "elfte|NUM": "5", "schack|NOUN": "5", "benägenhet|NOUN": "5", "intag|NOUN": "5", "stadion|NOUN": "5", "autentisk|ADJ": "5", "blankett|NOUN": "5", "fotografering|NOUN": "5", "rullstol|NOUN": "5", "årtal|NOUN": "5", "språng|NOUN": "5", "brunn|NOUN": "5", "artificiell|ADJ": "5", "företagsamhet|NOUN": "5", "filtrera|VERB": "5", "förolämpning|NOUN": "5", "kompani|NOUN": "6", "subventionera|VERB": "5", "uthållighet|NOUN": "5", "matsal|NOUN": "5", "skymning|NOUN": "5", "bekvämlighet|NOUN": "5", "eländig|ADJ": "5", "ark|NOUN": "6", "bulle|NOUN": "5", "parad|NOUN": "5", "stressa|VERB": "5", "glimt|NOUN": "5", "massaker|NOUN": "5", "riklig|ADJ": "5", "utlopp|NOUN": "5", "diplomati|NOUN": "5", "sås|NOUN": "5", "omfamna|VERB": "5", "absorbera|VERB": "5", "brandman|NOUN": "5", "lätthet|NOUN": "5", "uppslutning|NOUN": "5", "farväl|NOUN": "5", "specificera|VERB": "5", "broms|NOUN": "5", "dynasti|NOUN": "5", "tomrum|NOUN": "5", "förbrukning|NOUN": "5", "klia|VERB": "5", "tillgripa|VERB": "5", "trög|ADJ": "5", "välgörenhet|NOUN": "5", "instinkt|NOUN": "5", "hädanefter|ADV": "5", "utdela|VERB": "5", "adoption|NOUN": "5", "försvinnande|NOUN": "5", "gisslan|NOUN": "5", "kvalificera|VERB": "5", "nykomling|NOUN": "5", "prenumeration|NOUN": "5", "barack|NOUN": "5", "fotbollsspelare|NOUN": "5", "förevändning|NOUN": "5", "aha|INTJ": "5", "bukt|NOUN": "5", "grundtanke|NOUN": "5", "slicka|VERB": "5", "genial|ADJ": "5", "grind|NOUN": "5", "kuvert|NOUN": "5", "odödlig|ADJ": "5", "elektronik|NOUN": "5", "publicitet|NOUN": "5", "barnmorska|NOUN": "5", "påfallande|ADJ": "5", "kavaj|NOUN": "5", "lins|NOUN": "5", "psyke|NOUN": "5", "allergi|NOUN": "5", "resande|ADJ": "5", "specialisera|VERB": "5", "mognad|NOUN": "5", "skelett|NOUN": "5", "mager|ADJ": "5", "beslutsamhet|NOUN": "5", "brödraskap|NOUN": "5", "slumpmässig|ADJ": "5", "helgdag|NOUN": "5", "inlärning|NOUN": "5", "manuskript|NOUN": "5", "massvis|ADV": "5", "uppvisning|NOUN": "5", "följeslagare|NOUN": "5", "ovetande|ADJ": "5", "portfölj|NOUN": "5", "trohet|NOUN": "5", "kontant|ADJ": "5", "kontanter|NOUN": "5", "bomull|NOUN": "5", "höna|NOUN": "5", "nattvard|NOUN": "5", "rutt|NOUN": "5", "avsättning|NOUN": "5", "lår|NOUN": "5", "motbevisa|VERB": "5", "gröt|NOUN": "5", "logotyp|NOUN": "5", "nyårsafton|NOUN": "5", "fläkt|NOUN": "5", "högtalare|NOUN": "5", "kräkas|VERB": "5", "lokalisera|VERB": "5", "lantbruk|NOUN": "5", "fjäril|NOUN": "5", "officer|NOUN": "5", "påbud|NOUN": "5", "underkläder|NOUN": "5", "hastig|ADJ": "5", "faster|NOUN": "5", "sammankalla|VERB": "5", "anekdot|NOUN": "5", "rekommenderad|ADJ": "5", "dike|NOUN": "5", "parfym|NOUN": "5", "intuition|NOUN": "5", "kortvarig|ADJ": "5", "växthus|NOUN": "5", "modul|NOUN": "5", "fantisera|VERB": "5", "landsman|NOUN": "5", "skönlitteratur|NOUN": "5", "maka|NOUN": "5", "prosa|NOUN": "5", "användbarhet|NOUN": "5", "förläggare|NOUN": "5", "förolämpa|VERB": "5", "påföljande|ADJ": "5", "notering|NOUN": "5", "nål|NOUN": "5", "talrik|ADJ": "5", "komplettering|NOUN": "5", "ordspråk|NOUN": "5", "solnedgång|NOUN": "5", "attribut|NOUN": "5", "fosterland|NOUN": "5", "klot|NOUN": "5", "utbetala|VERB": "5", "alfabet|NOUN": "5", "bokföring|NOUN": "5", "fräck|ADJ": "5", "gammaldags|ADJ": "5", "Jorden|PROPN": "5", "jaså|INTJ": "5", "lämplighet|NOUN": "5", "sönderfall|NOUN": "5", "ämbetsman|NOUN": "5", "duell|NOUN": "5", "likviditet|NOUN": "5", "lossna|VERB": "5", "mikrofon|NOUN": "5", "trottoar|NOUN": "5", "slips|NOUN": "5", "hormon|NOUN": "5", "illamående|NOUN": "5", "tilldelning|NOUN": "5", "aluminium|NOUN": "5", "kappa|NOUN": "5", "permission|NOUN": "5", "försprång|NOUN": "5", "intim|ADJ": "5", "älskare|NOUN": "5", "skvaller|NOUN": "5", "metodik|NOUN": "5", "attraktion|NOUN": "5", "fragment|NOUN": "5", "magister|NOUN": "5", "reserv|NOUN": "5", "ekologi|NOUN": "5", "sponsring|NOUN": "5", "adelsman|NOUN": "5", "maskineri|NOUN": "5", "spalt|NOUN": "5", "underkastelse|NOUN": "5", "uråldrig|ADJ": "5", "clown|NOUN": "5", "noll|NOUN": "5", "verbal|ADJ": "5", "framträdande|NOUN": "5", "polisstation|NOUN": "5", "borsta|VERB": "5", "bägare|NOUN": "5", "gränslös|ADJ": "5", "kärl|NOUN": "5", "utomordentlig|ADJ": "5", "manager|NOUN": "5", "sångerska|NOUN": "5", "kooperativ|NOUN": "5", "genomskinlig|ADJ": "5", "kalender|NOUN": "5", "option|NOUN": "5", "arkeolog|NOUN": "5", "oändlighet|NOUN": "5", "netto|NOUN": "5", "veto|NOUN": "5", "veteran|NOUN": "5", "kalori|NOUN": "5", "vits|NOUN": "5", "kruka|NOUN": "5", "lotteri|NOUN": "5", "spektrum|NOUN": "5", "attentat|NOUN": "5", "avtala|VERB": "5", "förutsägelse|NOUN": "5", "halvtid|NOUN": "5", "kvitto|NOUN": "5", "oförutsedd|ADJ": "5", "livskraftig|ADJ": "5", "delegera|VERB": "5", "flit|NOUN": "5", "fullvärdig|ADJ": "5", "stab|NOUN": "5", "päron|NOUN": "5", "myndig|ADJ": "5", "förräderi|NOUN": "5", "förskott|NOUN": "5", "raka|VERB": "5", "svida|VERB": "5", "syntetisk|ADJ": "5", "mala|VERB": "5", "frisör|NOUN": "5", "osanning|NOUN": "5", "identifiering|NOUN": "5", "undre|ADJ": "5", "återvinning|NOUN": "5", "hurra|VERB": "5", "landning|NOUN": "5", "spilla|VERB": "5", "duva|NOUN": "5", "pryda|VERB": "5", "karakterisera|VERB": "5", "komponera|VERB": "5", "vidsträckt|ADJ": "5", "areal|NOUN": "5", "utvecklare|NOUN": "5", "betjäna|VERB": "5", "projektion|NOUN": "5", "skrattretande|ADJ": "5", "bacon|NOUN": "5", "gräl|NOUN": "5", "diameter|NOUN": "5", "förhöra|VERB": "5", "läsk|NOUN": "5", "tillmäta|VERB": "5", "åsna|NOUN": "5", "konsolidering|NOUN": "5", "tidtabell|NOUN": "5", "återbetalning|NOUN": "5", "explicit|ADV": "5", "kafé (el. café)|NOUN": "5", "manifest|ADJ": "5", "stram|ADJ": "5", "handske|NOUN": "5", "informativ|ADJ": "5", "rekonstruktion|NOUN": "5", "ridning|NOUN": "5", "garn|NOUN": "5", "samtidig|ADJ": "5", "matt|ADJ": "5", "bredda|VERB": "5", "gruppledare|NOUN": "5", "certifikat|NOUN": "5", "garage|NOUN": "5", "sociologi|NOUN": "5", "angränsande|ADJ": "5", "festlig|ADJ": "5", "generalisera|VERB": "5", "glödlampa|NOUN": "5", "grubbla|VERB": "5", "lantbrukare|NOUN": "5", "stipendium|NOUN": "5", "strukturera|VERB": "5", "tjur|NOUN": "5", "böna|NOUN": "5", "erotisk|ADJ": "5", "förträfflig|ADJ": "5", "löpare|NOUN": "5", "medlidande|NOUN": "5", "spänd|ADJ": "5", "gardin|NOUN": "5", "programmerare|NOUN": "5", "radiostation|NOUN": "5", "hosta|VERB": "5", "jämvikt|NOUN": "5", "tonvikt|NOUN": "5", "lobby|NOUN": "5", "explosiv|ADJ": "5", "hjälplös|ADJ": "5", "klausul|NOUN": "5", "spindel|NOUN": "5", "topplista|NOUN": "5", "klump|NOUN": "5", "trivsam|ADJ": "5", "brådskande|ADJ": "5", "elementär|ADJ": "5", "rättfärdiga|VERB": "5", "navigera|VERB": "5", "darra|VERB": "5", "flygel|NOUN": "5", "orientering|NOUN": "5", "utpräglad|ADJ": "5", "bebo|VERB": "5", "embryo|NOUN": "5", "lexikon|NOUN": "5", "experimentell|ADJ": "5", "instifta|VERB": "5", "väsentligen|ADV": "5", "kortfattad|ADJ": "5", "referat|NOUN": "5", "fyr|NOUN": "5", "förbränning|NOUN": "5", "inrymma|VERB": "5", "privilegierad|ADJ": "5", "kardinal|NOUN": "5", "essens|NOUN": "5", "affärsverksamhet|NOUN": "5", "extraordinär|ADJ": "5", "grammatik|NOUN": "5", "komposition|NOUN": "5", "krok|NOUN": "5", "kyss|NOUN": "5", "företrädesvis|ADV": "5", "medfödd|ADJ": "5", "jurisdiktion|NOUN": "5", "knipa|VERB": "5", "kondition|NOUN": "5", "oriktig|ADJ": "5", "proportionell|ADJ": "5", "själslig|ADJ": "5", "dagsljus|NOUN": "5", "fukt|NOUN": "5", "abonnemang|NOUN": "5", "sammanföra|VERB": "5", "ånga|NOUN": "5", "aktiemarknad|NOUN": "5", "mapp|NOUN": "5", "prototyp|NOUN": "5", "vilseleda|VERB": "5", "immigrant|NOUN": "5", "anlag|NOUN": "5", "fullmakt|NOUN": "5", "hyresvärd|NOUN": "5", "klassificering|NOUN": "5", "parlamentsledamot|NOUN": "5", "försena|VERB": "5", "renhet|NOUN": "5", "övertid|NOUN": "6", "allergisk|ADJ": "6", "eskalera|VERB": "6", "föreståndare|NOUN": "6", "spanare|NOUN": "6", "instruktör|NOUN": "6", "mugg|NOUN": "6", "granat|NOUN": "6", "ofrivillig|ADJ": "6", "subtil|ADJ": "6", "successiv|ADJ": "6", "välvilja|NOUN": "6", "banal|ADJ": "6", "spjut|NOUN": "6", "hektar|NOUN": "6", "avvärja|VERB": "6", "hållplats|NOUN": "6", "härma|VERB": "6", "distributör|NOUN": "6", "hårdvara|NOUN": "6", "grop|NOUN": "6", "repetera|VERB": "6", "utrotning|NOUN": "6", "grannskap|NOUN": "6", "kamel|NOUN": "6", "avlopp|NOUN": "6", "hjälpsam|ADJ": "6", "ämnesområde|NOUN": "6", "ändlös|ADJ": "6", "flamma|NOUN": "6", "livmoder|NOUN": "6", "reduktion|NOUN": "6", "susa|VERB": "6", "funktionalitet|NOUN": "6", "kulminera|VERB": "6", "slät|ADJ": "6", "hysteri|NOUN": "6", "rulle|NOUN": "6", "nattlig|ADJ": "6", "stråle|NOUN": "6", "avskilja|VERB": "6", "värdesätta|VERB": "6", "bark|NOUN": "6", "nalle|NOUN": "6", "fångst|NOUN": "6", "revolutionerande|ADJ": "6", "fåtölj|NOUN": "6", "ogiltig|ADJ": "6", "hygien|NOUN": "6", "tegel|NOUN": "6", "accelerera|VERB": "6", "gedigen|ADJ": "6", "känslighet|NOUN": "6", "sluttning|NOUN": "6", "nordväst|NOUN": "6", "utsökt|ADJ": "6", "analogi|NOUN": "6", "specifikation|NOUN": "6", "samordnare|NOUN": "6", "stöt|NOUN": "6", "bandit|NOUN": "6", "devalvering|NOUN": "6", "internationalisering|NOUN": "6", "kölvatten|NOUN": "6", "frige|VERB": "6", "åska|NOUN": "6", "hallå|NOUN": "6", "badkar|NOUN": "6", "obligation|NOUN": "6", "vertikal|ADJ": "6", "sommarlov|NOUN": "6", "volontär|NOUN": "6", "likgiltighet|NOUN": "6", "mottaglig|ADJ": "6", "noggrannhet|NOUN": "6", "tjat|NOUN": "6", "addera|VERB": "6", "barnvagn|NOUN": "6", "hurra|INTJ": "6", "simning|NOUN": "6", "omvårdnad|NOUN": "6", "beskydda|VERB": "6", "fyrkantig|ADJ": "6", "tunna|NOUN": "6", "ull|NOUN": "6", "avresa|NOUN": "6", "båge|NOUN": "6", "robust|ADJ": "6", "suppleant|NOUN": "6", "energisk|ADJ": "6", "rikligt|ADV": "6", "blotta|VERB": "6", "lokalisering|NOUN": "6", "interagera|VERB": "6", "julgran|NOUN": "6", "porto|NOUN": "6", "stick|NOUN": "6", "rotera|VERB": "6", "kiosk|NOUN": "6", "galler|NOUN": "6", "onormal|ADJ": "6", "oräknelig|ADJ": "6", "olivolja|NOUN": "6", "bokning|NOUN": "6", "förskräcklig|ADJ": "6", "inspektera|VERB": "6", "orientera|VERB": "6", "smeka|VERB": "6", "välgörande|ADJ": "6", "reception|NOUN": "6", "reproduktion|NOUN": "6", "konsul|NOUN": "6", "konsulat|NOUN": "6", "medvetslös|ADJ": "6", "moped|NOUN": "6", "sammanträda|VERB": "6", "altare|NOUN": "6", "kidnappning|NOUN": "6", "uppfyllelse|NOUN": "6", "betingelse|NOUN": "6", "förplikta|VERB": "6", "handväska|NOUN": "6", "häkta|VERB": "6", "rådjur|NOUN": "6", "specialisering|NOUN": "6", "överfall|NOUN": "6", "frimärke|NOUN": "6", "lakan|NOUN": "6", "gurka|NOUN": "6", "kanna|NOUN": "6", "midja|NOUN": "6", "omringa|VERB": "6", "styrelseordförande|NOUN": "6", "ödelägga|VERB": "6", "slang|NOUN": "6", "överhuvud|NOUN": "6", "handelsman|NOUN": "6", "linjär|ADJ": "6", "telekommunikation|NOUN": "6", "karakteristisk|ADJ": "6", "åklagarmyndighet|NOUN": "6", "årsdag|NOUN": "6", "repetition|NOUN": "6", "underskrift|NOUN": "6", "förgrund|NOUN": "6", "grönska|NOUN": "6", "kungörelse|NOUN": "6", "besvära|VERB": "6", "reflex|NOUN": "6", "inspektör|NOUN": "6", "stum|ADJ": "6", "uppdra|VERB": "6", "gunga|VERB": "6", "kooperativ|ADJ": "6", "legitimation|NOUN": "6", "patriotisk|ADJ": "6", "aptit|NOUN": "6", "artig|ADJ": "6", "beskyddare|NOUN": "6", "samstämmighet|NOUN": "6", "uppehälle|NOUN": "6", "segment|NOUN": "6", "stege|NOUN": "6", "rea|NOUN": "6", "oliv|NOUN": "6", "syra|NOUN": "6", "vattna|VERB": "6", "besätta|VERB": "6", "dispyt|NOUN": "6", "kräfta|NOUN": "6", "läcker|ADJ": "6", "vaktmästare|NOUN": "6", "byggnation|NOUN": "6", "förlåt|INTJ": "6", "bi|NOUN": "6", "dårskap|NOUN": "6", "räka|NOUN": "6", "terminal|NOUN": "6", "vakuum|NOUN": "6", "fusion|NOUN": "6", "utskrift|NOUN": "6", "offert|NOUN": "6", "botemedel|NOUN": "6", "säregen|ADJ": "6", "taxa|NOUN": "6", "välvillig|ADJ": "6", "klumpig|ADJ": "6", "tillflykt|NOUN": "6", "vävnad|NOUN": "6", "majestät|NOUN": "6", "immunitet|NOUN": "6", "ombildning|NOUN": "6", "omstridd|ADJ": "6", "periferi|NOUN": "6", "nunna|NOUN": "6", "löjtnant|NOUN": "6", "återlämna|VERB": "6", "stav|NOUN": "6", "fridfull|ADJ": "6", "höghus|NOUN": "6", "innevånare|NOUN": "6", "sjösätta|VERB": "6", "trauma|NOUN": "6", "oväder|NOUN": "6", "spion|NOUN": "6", "komplicera|VERB": "6", "substantiv|NOUN": "6", "undersida|NOUN": "6", "putsa|VERB": "6", "kam|NOUN": "6", "manuell|ADJ": "6", "mittfält|NOUN": "6", "pizzeria|NOUN": "6", "sittplats|NOUN": "6", "uthyrning|NOUN": "6", "komplimang|NOUN": "6", "handtag|NOUN": "6", "bemästra|VERB": "6", "obekant|ADJ": "6", "stapla|VERB": "6", "tusental|NOUN": "6", "berättiga|VERB": "6", "stereotyp|ADJ": "6", "vitlök|NOUN": "6", "alkoholism|NOUN": "6", "beröring|NOUN": "6", "bete|NOUN": "6", "flerårig|ADJ": "6", "förråda|VERB": "6", "försändelse|NOUN": "6", "resväska|NOUN": "6", "flyktig|ADJ": "6", "kirurg|NOUN": "6", "otvivelaktigt|ADV": "6", "saft|NOUN": "6", "varaktighet|NOUN": "6", "lekplats|NOUN": "6", "tillförlitlighet|NOUN": "6", "adjö|INTJ": "6", "käpp|NOUN": "6", "lossa|VERB": "6", "summering|NOUN": "6", "exekutiv|ADJ": "6", "kandidatur|NOUN": "6", "tum|NOUN": "6", "återkoppling|NOUN": "6", "dofta|VERB": "6", "encyklopedi|NOUN": "6", "förrädare|NOUN": "6", "tvättmaskin|NOUN": "6", "kvist|NOUN": "6", "tvål|NOUN": "6", "madrass|NOUN": "6", "heder|NOUN": "6", "knop|NOUN": "6", "maträtt|NOUN": "6", "njure|NOUN": "6", "alstra|VERB": "6", "beslutsam|ADJ": "6", "kontur|NOUN": "6", "värka|VERB": "6", "droppe|NOUN": "6", "inställa|VERB": "6", "programmera|VERB": "6", "resebyrå|NOUN": "6", "gnista|NOUN": "6", "envishet|NOUN": "6", "stilig|ADJ": "6", "vänskaplig|ADJ": "6", "kristall|NOUN": "6", "passionerad|ADJ": "6", "yr|ADJ": "6", "besiktning|NOUN": "6", "delgivning|NOUN": "6", "gjuta|VERB": "6", "smörja|VERB": "6", "ådra|VERB": "6", "åkomma|NOUN": "6", "stång|NOUN": "6", "konsultera|VERB": "6", "återuppliva|VERB": "6", "växtlighet|NOUN": "6", "frost|NOUN": "6", "lykta|NOUN": "6", "akustisk|ADJ": "6", "antydning|NOUN": "6", "häl|NOUN": "6", "hängivenhet|NOUN": "6", "orätt|NOUN": "6", "syntes|NOUN": "6", "ungdomlig|ADJ": "6", "citron|NOUN": "6", "tillbakadragande|NOUN": "6", "förfalskning|NOUN": "6", "tass|NOUN": "6", "trasa|NOUN": "6", "orgel|NOUN": "6", "oberoende|NOUN": "6", "geometri|NOUN": "6", "omfång|NOUN": "6", "oviss|ADJ": "6", "uteslutning|NOUN": "6", "utsända|VERB": "6", "pensionering|NOUN": "6", "förstora|VERB": "6", "försvinnande|ADV": "6", "paraply|NOUN": "6", "plakat|NOUN": "6", "veranda|NOUN": "6", "kosttillskott|NOUN": "6", "krock|NOUN": "6", "skyltfönster|NOUN": "6", "munter|ADJ": "6", "shorts|NOUN": "6", "vandrarhem|NOUN": "6", "kvadrat|NOUN": "6", "raseri|NOUN": "6", "tangent|NOUN": "6", "interiör|NOUN": "6", "bondgård|NOUN": "6", "brådska|NOUN": "6", "svartsjuka|NOUN": "6", "älskarinna|NOUN": "6", "adjektiv|NOUN": "6", "berömmelse|NOUN": "6", "bundsförvant|NOUN": "6", "fjärran|ADV": "6", "utantill|ADV": "6", "överträda|VERB": "6", "bortskämd|ADJ": "6", "byggare|NOUN": "6", "obildad|ADJ": "6", "bål|NOUN": "6", "horisontell|ADJ": "6", "imitera|VERB": "6", "optisk|ADJ": "6", "temperament|NOUN": "6", "uppställning|NOUN": "6", "bedragare|NOUN": "6", "tonfall|NOUN": "6", "fotografisk|ADJ": "6", "skissera|VERB": "6", "kollision|NOUN": "6", "magnetisk|ADJ": "6", "sparsam|ADJ": "6", "prestigefylld|ADJ": "6", "kran|NOUN": "6", "småstad|NOUN": "6", "vingård|NOUN": "6", "flamma|VERB": "6", "försona|VERB": "6", "treårig|ADJ": "6", "utlämna|VERB": "6", "linne|NOUN": "6", "nybyggare|NOUN": "6", "triangel|NOUN": "6", "utsliten|ADJ": "6", "slank|ADJ": "6", "annullera|VERB": "6", "brandkår|NOUN": "6", "pinne|NOUN": "6", "hare|NOUN": "6", "jämförande|ADJ": "6", "ministerium|NOUN": "6", "vikarie|NOUN": "6", "astma|NOUN": "6", "förvirra|VERB": "6", "inflammation|NOUN": "6", "larma|VERB": "6", "mätta|VERB": "6", "plåster|NOUN": "6", "rotation|NOUN": "6", "skolgård|NOUN": "6", "åtkomst|NOUN": "6", "övernatta|VERB": "6", "egenhet|NOUN": "6", "oordning|NOUN": "6", "revidering|NOUN": "6", "smörja|NOUN": "6", "ålderdom|NOUN": "6", "kommando|NOUN": "6", "utmattning|NOUN": "6", "keramik|NOUN": "6", "mustasch|NOUN": "6", "baron|NOUN": "6", "boss|NOUN": "6", "läder|NOUN": "6", "rengöring|NOUN": "6", "avfärd|NOUN": "6", "hink|NOUN": "6", "matematiker|NOUN": "6", "passning|NOUN": "6", "tillsättning|NOUN": "6", "hemort|NOUN": "6", "instruera|VERB": "6", "rengöra|VERB": "6", "dekoration|NOUN": "6", "månatlig|ADJ": "6", "patriotism|NOUN": "6", "tillmötesgå|VERB": "6", "gås|NOUN": "6", "programmering|NOUN": "6", "vicepresident|NOUN": "6", "avla|VERB": "6", "brigad|NOUN": "6", "allsidig|ADJ": "6", "komfort|NOUN": "6", "listig|ADJ": "6", "simulering|NOUN": "6", "återbetala|VERB": "6", "sned|ADJ": "6", "bassäng|NOUN": "6", "närbelägen|ADJ": "6", "pensel|NOUN": "6", "luftfart|NOUN": "6", "patrull|NOUN": "6", "arbetsrum|NOUN": "6", "implementering|NOUN": "6", "hydda|NOUN": "6", "oerfaren|ADJ": "6", "bokstavlig|ADJ": "6", "elektromagnetisk|ADJ": "6", "rymlig|ADJ": "6", "världsåskådning|NOUN": "6", "ansiktsuttryck|NOUN": "6", "frigivning|NOUN": "6", "pristagare|NOUN": "6", "självsäker|ADJ": "6", "fiber|NOUN": "6", "dricks|NOUN": "6", "tam|ADJ": "6", "oreda|NOUN": "6", "förnekande|NOUN": "6", "algoritm|NOUN": "6", "tall|NOUN": "6", "avsiktlig|ADJ": "6", "biolog|NOUN": "6", "tarm|NOUN": "6", "adlig|ADJ": "6", "spegelbild|NOUN": "6", "campus|NOUN": "6", "brännvin|NOUN": "6", "kompatibel|ADJ": "6", "ängslig|ADJ": "6", "tolfte|NUM": "6", "beväpna|VERB": "6", "tvåhundra|NUM": "6", "biff|NOUN": "6", "ratificering|NOUN": "6", "skådespelerska|NOUN": "6", "slavisk|ADJ": "6", "glänsa|VERB": "6", "ömhet|NOUN": "6", "föräldralös|ADJ": "6", "tumör|NOUN": "6", "vidareutveckling|NOUN": "6", "juice|NOUN": "6", "deponera|VERB": "6", "kirurgi|NOUN": "6", "närmande|NOUN": "6", "rondell|NOUN": "6", "sensationell|ADJ": "6", "stabilisering|NOUN": "6", "törst|NOUN": "6", "arkitektonisk|ADJ": "6", "förbluffande|ADV": "6", "klunga|NOUN": "6", "medfölja|VERB": "6", "processor|NOUN": "6", "tabu|ADJ": "6", "vulgär|ADJ": "6", "minnesmärke|NOUN": "6", "provision|NOUN": "6", "blödning|NOUN": "6", "defekt|NOUN": "6", "disposition|NOUN": "6", "koordinera|VERB": "6", "staket|NOUN": "6", "hytt|NOUN": "6", "kastrull|NOUN": "6", "startpunkt|NOUN": "6", "sked|NOUN": "6", "bal|NOUN": "6", "sandstrand|NOUN": "6", "stereotyp|NOUN": "6", "tålmodigt|ADV": "6", "arrestering|NOUN": "6", "kryssning|NOUN": "6", "pipa|VERB": "6", "gräla|VERB": "6", "area|NOUN": "6", "förbipasserande|ADJ": "6", "förlikning|NOUN": "6", "ljuda|VERB": "6", "samexistens|NOUN": "6", "terapeutisk|ADJ": "6", "trendig|ADJ": "6", "återhållsamhet|NOUN": "6", "hjort|NOUN": "6", "debitera|VERB": "6", "dundra|VERB": "6", "kräm|NOUN": "6", "korrespondent|NOUN": "6", "aktualitet|NOUN": "6", "behållare|NOUN": "6", "gruvarbetare|NOUN": "6", "åtstramning|NOUN": "6", "kontinental|ADJ": "6", "väster|NOUN": "6", "ankare|NOUN": "6", "åker|NOUN": "6", "senator|NOUN": "6", "häpnad|NOUN": "6", "mynning|NOUN": "6", "omtänksam|ADJ": "6", "omåttlig|ADJ": "6", "rekonstruera|VERB": "6", "maximum|NOUN": "6", "karaktärsdrag|NOUN": "6", "perfektion|NOUN": "6", "timmer|NOUN": "6", "urin|NOUN": "6", "arkivera|VERB": "6", "oavbruten|ADJ": "6", "kolonn|NOUN": "6", "appell|NOUN": "6", "strejka|VERB": "6", "propp|NOUN": "6", "automat|NOUN": "6", "studium|NOUN": "6", "högljudd|ADJ": "6", "skaldjur|NOUN": "6", "stinka|VERB": "6", "tillfreds|ADJ": "6", "världsomfattande|ADJ": "6", "befruktning|NOUN": "6", "glänsande|ADJ": "6", "organisatör|NOUN": "6", "pussel|NOUN": "6", "vitamin|NOUN": "6", "aktning|NOUN": "6", "boplats|NOUN": "6", "vederbörlig|ADJ": "6", "dråp|NOUN": "6", "jubileum|NOUN": "6", "frikänna|VERB": "6", "hetta|VERB": "6", "formation|NOUN": "6", "ridå|NOUN": "6", "rådfråga|VERB": "6", "svälla|VERB": "6", "avföring|NOUN": "6", "modifikation|NOUN": "6", "ordförråd|NOUN": "6", "tjocklek|NOUN": "6", "metropol|NOUN": "6", "injektion|NOUN": "6", "lantlig|ADJ": "6", "veckotidning|NOUN": "6", "orkester|NOUN": "6", "skruv|NOUN": "6", "solsken|NOUN": "6", "matvara|NOUN": "6", "regemente|NOUN": "6", "sammanträffande|NOUN": "6", "utstrålning|NOUN": "6", "valla|VERB": "6", "arvode|NOUN": "6", "periodisk|ADJ": "6", "favör|NOUN": "6", "kommunikativ|ADJ": "6", "terminal|ADJ": "6", "trappsteg|NOUN": "6", "paj|NOUN": "6", "anskaffa|VERB": "6", "mörkhyad|ADJ": "6", "tristess|NOUN": "6", "kassett|NOUN": "6", "räddare|NOUN": "6", "almanacka|NOUN": "6", "accent|NOUN": "6", "kvällsmat|NOUN": "6", "bestiga|VERB": "6", "styv|ADJ": "6", "knekt|NOUN": "6", "väv|NOUN": "6", "översvämma|VERB": "6", "örn|NOUN": "6", "seglare|NOUN": "6", "spöke|NOUN": "6", "lund|NOUN": "6", "tålmodig|ADJ": "6", "koja|NOUN": "6", "lockelse|NOUN": "6", "lärd|ADJ": "6", "balk|NOUN": "6", "åldring|NOUN": "6", "fullmåne|NOUN": "6", "bröstkorg|NOUN": "6", "slätt|ADV": "6", "spektakel|NOUN": "6", "ven|NOUN": "6", "nöt|NOUN": "6", "odjur|NOUN": "6", "äventyrare|NOUN": "6", "bildlig|ADJ": "6", "rangordna|VERB": "6", "smörgås|NOUN": "6", "hjord|NOUN": "6", "vildsvin|NOUN": "6", "bibliografi|NOUN": "6", "ihärdig|ADJ": "6", "indignation|NOUN": "6", "paradoxal|ADJ": "6", "soluppgång|NOUN": "6", "grädda|VERB": "6", "kontrovers|NOUN": "6", "multiplicera|VERB": "6", "oförrätt|NOUN": "6", "revben|NOUN": "6", "yoghurt|NOUN": "6", "delikat|ADJ": "6", "konsultation|NOUN": "6", "kväve|NOUN": "6", "kvarn|NOUN": "6", "gummi|NOUN": "6", "facilitet|NOUN": "6", "mittemot (el. mitt emot)|ADP": "6", "oenig|ADJ": "6", "oföränderlig|ADJ": "6", "restaurering|NOUN": "6", "snuskig|ADJ": "6", "tågstation|NOUN": "6", "herde|NOUN": "6", "kål|NOUN": "6", "tillförsel|NOUN": "6", "avskrivning|NOUN": "6", "bemanning|NOUN": "6", "pytteliten|ADJ": "6", "cirkulation|NOUN": "6", "termisk|ADJ": "6", "ömtålig|ADJ": "6", "koda|VERB": "6", "kämpe|NOUN": "6", "besatthet|NOUN": "6", "fjärrkontroll|NOUN": "6", "juvel|NOUN": "6", "ponny|NOUN": "6", "bemanna|VERB": "6", "måtta|NOUN": "6", "dekorera|VERB": "6", "gaffel|NOUN": "6", "pilgrim|NOUN": "6", "ackumulera|VERB": "6", "getto|NOUN": "6", "skorsten|NOUN": "6", "antenn|NOUN": "6", "montering|NOUN": "6", "synbar|ADJ": "6", "vrå|NOUN": "6", "assistera|VERB": "6", "defensiv|NOUN": "6", "videokamera|NOUN": "6", "bataljon|NOUN": "6", "intelligens|NOUN": "6", "diplom|NOUN": "6", "konfiguration|NOUN": "6", "efterfölja|VERB": "6", "exemplarisk|ADJ": "6", "konsistens|NOUN": "6", "stelna|VERB": "6", "amortering|NOUN": "6", "avskrift|NOUN": "6", "bläck|NOUN": "6", "restaurera|VERB": "6", "pulver|NOUN": "6", "remsa|NOUN": "6", "apelsin|NOUN": "6", "cement|NOUN": "6", "trailer|NOUN": "6", "ljum|ADJ": "6", "sammanstötning|NOUN": "6", "stormig|ADJ": "6", "pina|NOUN": "6", "skift|NOUN": "6", "stöna|VERB": "6", "uppsyn|NOUN": "6", "återse|VERB": "6", "elektron|NOUN": "6", "oanvändbar|ADJ": "6", "sömnig|ADJ": "6", "emission|NOUN": "6", "omloppsbana|NOUN": "6", "blixtsnabbt|ADV": "6", "brevväxling|NOUN": "6", "ventil|NOUN": "6", "fresta|VERB": "6", "pekfinger|NOUN": "6", "sigill|NOUN": "6", "armbåge|NOUN": "6", "ljusblå|ADJ": "6", "skaft|NOUN": "6", "paviljong|NOUN": "6", "segerrik|ADJ": "6", "skenbar|ADJ": "6", "svartsjuk|ADJ": "6", "mångfaldig|ADJ": "6", "omlopp|NOUN": "6", "kemist|NOUN": "6", "dykning|NOUN": "6", "orörlig|ADJ": "6", "tagning|NOUN": "6", "cykelväg|NOUN": "6", "donator|NOUN": "6", "förverkligande|NOUN": "6", "nyck|NOUN": "6", "gränsområde|NOUN": "6", "pittoresk|ADJ": "6", "yla|VERB": "6", "disciplinär|ADJ": "6", "farväl|INTJ": "6", "pånyttfödelse|NOUN": "6", "relik|NOUN": "6", "berättigande|NOUN": "6", "föresats|NOUN": "6", "inbetalning|NOUN": "6", "ströva|VERB": "6", "substitut|NOUN": "6", "tjugonde|NUM": "6", "arbetslag|NOUN": "6", "lim|NOUN": "6", "läglig|ADJ": "6", "nyttighet|NOUN": "6", "simhall|NOUN": "6", "animation|NOUN": "6", "väte|NOUN": "6", "orätt|ADJ": "6", "uppskov|NOUN": "6", "belägenhet|NOUN": "6", "sammandrag|NOUN": "6", "bensinstation|NOUN": "6", "gymnastik|NOUN": "6", "kommissarie|NOUN": "6", "vokal|NOUN": "6", "förmyndare|NOUN": "6", "mineral|NOUN": "6", "omnämnande|NOUN": "6", "alarm|NOUN": "6", "allé|NOUN": "6", "bergstopp|NOUN": "6", "navigation|NOUN": "6", "set|NOUN": "6", "tematisk|ADJ": "6", "täthet|NOUN": "6", "återupptäcka|VERB": "6", "postkontor|NOUN": "6", "ärm|NOUN": "6", "residens|NOUN": "6", "teleskop|NOUN": "6", "tryckning|NOUN": "6", "drickande|NOUN": "6", "kabinett|NOUN": "6", "charmerande|ADJ": "6", "missfall|NOUN": "6", "äktenskaplig|ADJ": "6", "emigrant|NOUN": "6", "bagatell|NOUN": "6", "bestämdhet|NOUN": "6", "aveny|NOUN": "6", "hosta|NOUN": "6", "andedräkt|NOUN": "6", "bottenvåning|NOUN": "6", "förtrolig|ADJ": "6", "avskedande|NOUN": "6", "femtonde|NUM": "6", "avbetalning|NOUN": "6", "fotgängare|NOUN": "6", "lärarinna|NOUN": "6", "terrass|NOUN": "6", "monter|NOUN": "6", "sylt|NOUN": "6", "kila|VERB": "6", "tuggummi|NOUN": "6", "bildskärm|NOUN": "6", "eliminering|NOUN": "6", "kalkylera|VERB": "6", "agentur|NOUN": "6", "mellanliggande|ADJ": "6", "trosa|NOUN": "6", "såg|NOUN": "6", "fysiologisk|ADJ": "6", "uppfödning|NOUN": "6", "betinga|VERB": "6", "farförälder|NOUN": "6", "råolja|NOUN": "6", "ficklampa|NOUN": "6", "hårig|ADJ": "6", "tvättmedel|NOUN": "6", "förorena|VERB": "6", "marskalk|NOUN": "6", "böjning|NOUN": "6", "narkoman|NOUN": "6", "upphetsning|NOUN": "6", "uppköp|NOUN": "6", "mentor|NOUN": "6", "fyrverkeri|NOUN": "6", "kollegium|NOUN": "6", "spade|NOUN": "6", "differentiering|NOUN": "6", "infektera|VERB": "6", "veck|NOUN": "6", "limma|VERB": "6", "oväsen|NOUN": "6", "innesluta|VERB": "6", "klädesplagg|NOUN": "6", "musiker|NOUN": "6", "smaklös|ADJ": "6", "stigning|NOUN": "6", "bravo|INTJ": "6", "hjärtlig|ADJ": "6", "explicit|ADJ": "6", "idrottsman|NOUN": "6", "koncession|NOUN": "6", "ofördelaktig|ADJ": "6", "ädel|ADJ": "6", "epos|NOUN": "6", "fasta|NOUN": "6", "geting|NOUN": "6", "hedervärd|ADJ": "6", "hjältinna|NOUN": "6", "knipa|NOUN": "6", "frågeformulär|NOUN": "6", "densitet|NOUN": "6", "eskortera|VERB": "6", "rankning|NOUN": "6", "servitör|NOUN": "6", "svägerska|NOUN": "6", "förbrylla|VERB": "6", "skattemässig|ADJ": "6", "tillgivenhet|NOUN": "6", "avkomling|NOUN": "6", "diagnostisera|VERB": "6", "rådman|NOUN": "6", "sammanfoga|VERB": "6", "ögonkast|NOUN": "6", "designer|NOUN": "6", "basilika|NOUN": "6", "lem|NOUN": "6", "adressera|VERB": "6", "bagare|NOUN": "6", "veckoslut|NOUN": "6", "centrera|VERB": "6", "fotfolk|NOUN": "6", "fästmö|NOUN": "6", "illvilja|NOUN": "6", "inskrivning|NOUN": "6", "omkrets|NOUN": "6", "självdeklaration|NOUN": "6", "trehundra|NUM": "6", "logo|NOUN": "6", "fyndighet|NOUN": "6", "gästfrihet|NOUN": "6", "konfirmation|NOUN": "6", "skär|NOUN": "6", "vindruva|NOUN": "6", "vårdare|NOUN": "6", "ådra|NOUN": "6", "tillfredsställd|ADJ": "6", "förestå|VERB": "6", "handflata|NOUN": "6", "inbillning|NOUN": "6", "logg|NOUN": "6", "bakverk|NOUN": "6", "gratulation|NOUN": "6", "kapplöpning|NOUN": "6", "opponent|NOUN": "6", "betydlig|ADJ": "6", "matris|NOUN": "6", "avdela|VERB": "6", "huvudämne|NOUN": "6", "komplott|NOUN": "6", "returnera|VERB": "6", "stadfästa|VERB": "6", "oavgjord|ADJ": "6", "beslutsamt|ADV": "6", "kupong|NOUN": "6", "massera|VERB": "6", "tändsticka|NOUN": "6", "ädelsten|NOUN": "6", "kakao|NOUN": "6", "akvarium|NOUN": "6", "smycke|NOUN": "6", "försvarsadvokat|NOUN": "6", "knytnäve|NOUN": "6", "optik|NOUN": "6", "skolkamrat|NOUN": "6", "synfält|NOUN": "6", "underlydande|ADJ": "6", "frist|NOUN": "6", "fyllning|NOUN": "6", "förvarna|VERB": "6", "stearinljus|NOUN": "6", "enhällig|ADJ": "6", "insjö|NOUN": "6", "ledsaga|VERB": "6", "moderskap|NOUN": "6", "undantagslöst|ADV": "6", "alldaglig|ADJ": "6", "avslappning|NOUN": "6", "konduktör|NOUN": "6", "lågstadium|NOUN": "6", "sportig|ADJ": "6", "utsändning|NOUN": "6", "villighet|NOUN": "6", "glans|NOUN": "6", "arvinge|NOUN": "6", "häfte|NOUN": "6", "mejeri|NOUN": "6", "chockera|VERB": "6", "eskort|NOUN": "6", "tabu|NOUN": "6", "avdelningschef|NOUN": "6", "pilgrimsfärd|NOUN": "6", "rättfram|ADJ": "6", "slaktare|NOUN": "6", "betecknande|ADJ": "6", "patologisk|ADJ": "6", "multimedia|NOUN": "6", "frånskild|ADJ": "6", "krämpa|NOUN": "6", "långsamhet|NOUN": "6", "mätare|NOUN": "6", "oljud|NOUN": "6", "slitage|NOUN": "6", "kommendant|NOUN": "6", "hök|NOUN": "6", "rugby|NOUN": "6", "snöre|NOUN": "6", "vidröra|VERB": "6", "dån|NOUN": "6", "sanitär|ADJ": "6", "stekpanna|NOUN": "6", "idol|NOUN": "6", "luftkonditionering|NOUN": "6", "svärson|NOUN": "6", "tejp|NOUN": "6", "viskning|NOUN": "6", "fatal|ADJ": "6", "arbetsam|ADJ": "6", "korporativ|ADJ": "6", "långfristig|ADJ": "6", "snarka|VERB": "6", "tunna|VERB": "6", "ärta|NOUN": "6", "kassaskåp|NOUN": "6", "fela|VERB": "6", "maskulin|ADJ": "6", "radie|NOUN": "6", "utväxling|NOUN": "6", "växellåda|NOUN": "6", "ånga|VERB": "6", "försyn|NOUN": "6", "glidning|NOUN": "6", "planlägga|VERB": "6", "feminin|ADJ": "6", "kodifiera|VERB": "6", "poem|NOUN": "6", "kompanjon|NOUN": "6", "stygg|ADJ": "6", "anstöt|NOUN": "6", "betyg(s)sätta|VERB": "6", "defekt|ADJ": "6", "fadd|ADJ": "6", "sittning|NOUN": "6", "besk|ADJ": "6", "rigorös|ADJ": "6", "moster|NOUN": "6", "gnida|VERB": "6", "ordningsföljd|NOUN": "6", "ärorik|ADJ": "6", "gnistra|VERB": "6", "pyjamas|NOUN": "6", "bergig|ADJ": "6", "fuktighet|NOUN": "6", "inkassera|VERB": "6", "laglighet|NOUN": "6", "statist|NOUN": "6", "nobel|ADJ": "6", "beväpning|NOUN": "6", "gymnasist|NOUN": "6", "kolossal|ADJ": "6", "stek|NOUN": "6", "uppkalla|VERB": "6", "försegla|VERB": "6", "konsortium|NOUN": "6", "acceptans|NOUN": "6", "grammatisk|ADJ": "6", "strykning|NOUN": "6", "kalcium|NOUN": "6", "fasta|VERB": "6", "tillfälligtvis|ADV": "6", "genomgående|ADV": "6", "hänförelse|NOUN": "6", "spårning|NOUN": "6", "systerson|NOUN": "6", "gunga|NOUN": "6", "ohyra|NOUN": "6", "opublicerad|ADJ": "6", "idrottsplats|NOUN": "6", "elastisk|ADJ": "6", "arrest|NOUN": "6", "dill|NOUN": "6", "vax|NOUN": "6", "pose|NOUN": "6", "bullrig|ADJ": "6", "spröd|ADJ": "6", "tidsskrift|NOUN": "6", "handfat|NOUN": "6", "kork|NOUN": "6", "immun|ADJ": "6", "inlämna|VERB": "6", "projektering|NOUN": "6", "regelbundenhet|NOUN": "6", "karavan|NOUN": "6", "krabba|NOUN": "6", "membran|NOUN": "6", "antikvitet|NOUN": "6", "brant|NOUN": "6", "genomträngande|ADJ": "6", "kemikalie|NOUN": "6", "kultiverad|ADJ": "6", "rumslig|ADJ": "6", "tråkighet|NOUN": "6", "namnteckning|NOUN": "6", "personell|ADJ": "6", "ungkarl|NOUN": "6", "rättfärdigande|NOUN": "6", "sammankoppla|VERB": "6", "aktivering|NOUN": "6", "mellantid|NOUN": "6", "motorbåt|NOUN": "6", "reglemente|NOUN": "6", "decimal|NOUN": "6", "mosa|VERB": "6", "olivträd|NOUN": "6", "anskaffning|NOUN": "6", "gradera|VERB": "6", "huva|NOUN": "6", "lodrät|ADJ": "6", "brodera|VERB": "6", "socka|NOUN": "6", "systerdotter|NOUN": "6", "turkos|NOUN": "6", "huvudrollsinnehavare|NOUN": "6", "kraftlös|ADJ": "6", "spann|NOUN": "6", "förbittring|NOUN": "6", "metallisk|ADJ": "6", "repertoar|NOUN": "6", "avspänd|ADJ": "6", "butiksägare|NOUN": "6", "kännare|NOUN": "6", "samtalspartner|NOUN": "6", "överväldiga|VERB": "6", "rea|VERB": "6", "böna|VERB": "6", "diagnostisk|ADJ": "6", "ställ|NOUN": "6", "kontingent|NOUN": "6", "projektil|NOUN": "6", "avtäcka|VERB": "6", "iakttagare|NOUN": "6", "atmosfärisk|ADJ": "6", "borttagning|NOUN": "6", "differentiera|VERB": "6", "fysiker|NOUN": "6", "mygga|NOUN": "6", "orange|NOUN": "6", "silke|NOUN": "6", "troende|NOUN": "6", "borste|NOUN": "6", "sparv|NOUN": "6", "stränghet|NOUN": "6", "nittonde|NUM": "6", "i övermorgon|ADV": "6", "motsägande|ADJ": "6", "käring|NOUN": "6", "blus|NOUN": "6", "kärnpunkt|NOUN": "6", "projektera|VERB": "6", "utstyrsel|NOUN": "6", "laser|NOUN": "6", "knippe|NOUN": "6", "presidium|NOUN": "6", "kvast|NOUN": "6", "plommon|NOUN": "6", "ägarskap|NOUN": "6", "oxe|NOUN": "6", "snabbköp|NOUN": "6", "tilltugg|NOUN": "6", "sned|NOUN": "6", "egenartad|ADJ": "6", "bulletin|NOUN": "6", "högerhand|NOUN": "6", "squash|NOUN": "6", "stadsbo|NOUN": "6", "simmare|NOUN": "6", "inkvartering|NOUN": "6", "majs|NOUN": "6", "visare|NOUN": "6", "oupphörlig|ADJ": "6", "bönfalla|VERB": "6", "dosering|NOUN": "6", "studiekamrat|NOUN": "6", "tryne|NOUN": "6", "ånger|NOUN": "6", "kvarlåtenskap|NOUN": "6", "körsbär|NOUN": "6", "rakning|NOUN": "6", "integral|NOUN": "6", "klibba|VERB": "6", "sparsamhet|NOUN": "6", "tunnland|NOUN": "6", "formge|VERB": "6", "moderlig|ADJ": "6", "pina|VERB": "6", "undervärdera|VERB": "6", "jetplan|NOUN": "6", "auktorisera|VERB": "6", "korporation|NOUN": "6", "saliv|NOUN": "6", "strömbrytare|NOUN": "6", "kurera|VERB": "6", "legering|NOUN": "6", "smaklig|ADJ": "6", "terroristisk|ADJ": "6", "hemgift|NOUN": "6", "avvara|VERB": "6", "förhandsvisning|NOUN": "6", "marmelad|NOUN": "6", "trafikpolis|NOUN": "6", "kittel|NOUN": "6", "bi|ADV": "6", "brådska|VERB": "6", "reseledare|NOUN": "6", "akustik|NOUN": "6", "forcerad|ADJ": "6", "tidsschema|NOUN": "6", "årtusende|NOUN": "6", "anträffa|VERB": "6", "rutnät|NOUN": "6", "försakelse|NOUN": "6", "pluton|NOUN": "6", "ägarinna|NOUN": "6", "överräcka|VERB": "6", "jordgubbe|NOUN": "6", "sesam|NOUN": "6", "artikulera|VERB": "6", "aprikos|NOUN": "6", "krage|NOUN": "6", "reklamera|VERB": "6", "tempus|NOUN": "6", "upplag|NOUN": "6", "tekniker|NOUN": "6", "avläsning|NOUN": "6", "knall|NOUN": "6", "molnig|ADJ": "6", "sårande|ADJ": "6", "särprägel|NOUN": "6", "variabel|ADJ": "6", "yrkesman|NOUN": "6", "återuppståndelse|NOUN": "6", "manöver|NOUN": "6", "myr|NOUN": "6", "överse|VERB": "6", "atletisk|ADJ": "6", "skolflicka|NOUN": "6", "atlet|NOUN": "6", "debitering|NOUN": "6", "huslig|ADJ": "6", "postlåda|NOUN": "6", "millennium|NOUN": "6", "valla|NOUN": "6", "armbandsur|NOUN": "6", "betäckning|NOUN": "6", "brorsdotter|NOUN": "6", "brutto|ADV": "6", "scarf|NOUN": "6", "annullering|NOUN": "6", "flanera|VERB": "6", "läkarvetenskap|NOUN": "6", "mittemot (el. mitt emot)|ADV": "6", "apparatur|NOUN": "6", "fosterbarn|NOUN": "6", "förbluffa|VERB": "6", "illamående|ADJ": "6", "vrist|NOUN": "6", "avskedsansökan|NOUN": "6", "blyertspenna|NOUN": "6", "invändig|ADJ": "6", "postulat|NOUN": "6", "ytterlig|ADJ": "6", "ungdomstid|NOUN": "6", "kabin|NOUN": "6", "nödhjälp|NOUN": "6", "kuriositet|NOUN": "6", "pantsätta|VERB": "6", "hake|NOUN": "6", "renlighet|NOUN": "6", "stjälk|NOUN": "6", "överlämning|NOUN": "6", "olympiad|NOUN": "6", "bräde|NOUN": "6", "hålighet|NOUN": "6", "realisering|NOUN": "6", "tariff|NOUN": "6", "bindel|NOUN": "6", "sockel|NOUN": "6", "animering|NOUN": "6", "didaktisk|ADJ": "6", "doktorsgrad|NOUN": "6", "husgeråd|NOUN": "6", "klarvaken|ADJ": "6", "bullra|VERB": "6", "persika|NOUN": "6", "svärdotter|NOUN": "6", "upprepat|ADV": "6", "genomskinlighet|NOUN": "6", "sonson|NOUN": "6", "stridslysten|ADJ": "6", "teatralisk|ADJ": "6", "tyngdkraft|NOUN": "6", "progression|NOUN": "6", "stadgande|NOUN": "6", "infarkt|NOUN": "6", "upphängning|NOUN": "6", "tesked|NOUN": "6", "uppdykande|ADJ": "6", "måtta|VERB": "6", "singularis|NOUN": "6", "dotterdotter|NOUN": "6", "syskonbarn|NOUN": "6", "veterinär|ADJ": "6", "baktala|VERB": "6", "påskrift|NOUN": "6", "slutta|VERB": "6", "farmaceutisk|ADJ": "6", "innertak|NOUN": "6", "knackning|NOUN": "6", "koffert|NOUN": "6", "monitor|NOUN": "6", "simbassäng|NOUN": "6", "trettionde|NUM": "6", "utvändig|ADJ": "6", "brudgum|NOUN": "6", "inneslutning|NOUN": "6", "genomresa|NOUN": "6", "karakteristik|NOUN": "6", "mör|ADJ": "6", "genomfart|NOUN": "6", "kameraman|NOUN": "6", "dotterson|NOUN": "6", "koefficient|NOUN": "6", "vägavgift|NOUN": "6", "adjö|NOUN": "6", "betjäning|NOUN": "6", "periodiskt|ADV": "6", "trofé|NOUN": "6", "vokal|ADJ": "6", "fjäder|NOUN": "6", "himmelsblå|ADJ": "6", "trådbuss|NOUN": "6", "trasa|VERB": "6", "födelsemärke|NOUN": "6", "hövlighet|NOUN": "6", "konvergens|NOUN": "6", "sorgsenhet|NOUN": "6", "brorson|NOUN": "6", "ringklocka|NOUN": "6", "vardaglighet|NOUN": "6", "berömdhet|NOUN": "6", "förutbestämma|VERB": "6", "folie|NOUN": "6", "kejsardöme|NOUN": "6", "käke|NOUN": "6", "rymling|NOUN": "6", "serum|NOUN": "6", "avresa|VERB": "6", "elektriker|NOUN": "6", "syrsa|NOUN": "6", "turkos|ADJ": "6", "äggvita|NOUN": "6", "hypotekslån|NOUN": "6", "invalid|NOUN": "6", "månljus|NOUN": "6", "transplantera|VERB": "6", "tursam|ADJ": "6", "kvalificering|NOUN": "6", "skolväska|NOUN": "6", "utprovning|NOUN": "6", "skollov|NOUN": "6", "likkista|NOUN": "6", "packe|NOUN": "6", "svärmor|NOUN": "6", "bäcken|NOUN": "6", "förbrukare|NOUN": "6", "grönska|VERB": "6", "modus|NOUN": "6", "studenthem|NOUN": "6", "mekaniker|NOUN": "6", "översida|NOUN": "6", "fullbordande|NOUN": "6", "undervåning|NOUN": "6", "aritmetisk|ADJ": "6", "fela|NOUN": "6", "frisersalong|NOUN": "6", "fönsterbräda|NOUN": "6", "cirkelformad|ADJ": "6", "kardinal|ADJ": "6", "oföränderligt|ADV": "6", "regelvidrig|ADJ": "6", "skrynkla|VERB": "6", "otvivelaktig|ADJ": "6", "sondotter|NOUN": "6", "ekolog|NOUN": "6", "åska|VERB": "6", "femtionde|NUM": "6", "gravera|VERB": "6", "ortopedi|NOUN": "6", "tekanna|NOUN": "6", "fyrtionde|NUM": "6", "konservator|NOUN": "6", "hurra|NOUN": "6", "inrikes|ADV": "6", "maka|VERB": "6", "askkopp|NOUN": "6", "fästman|NOUN": "6", "hyvel|NOUN": "6", "straffspark|NOUN": "6", "stött|ADJ": "6", "subtrahera|VERB": "6", "kakelplatta|NOUN": "6", "kasus|NOUN": "6", "svärfar|NOUN": "6", "dossier|NOUN": "6", "nolla|VERB": "6", "återgälda|VERB": "6", "besk|NOUN": "6", "bräda|VERB": "6", "dyrkan|NOUN": "6", "enfamiljshus|NOUN": "6", "förkroppsligande|NOUN": "6", "violin|NOUN": "6", "mottaga|VERB": "6", "nittionde|NUM": "6", "oregelbundenhet|NOUN": "6", "sjukskötare|NOUN": "6", "stockning|NOUN": "6", "toffel|NOUN": "6", "vattenmelon|NOUN": "6", "verkställare|NOUN": "6", "vårlig|ADJ": "6", "metalltråd|NOUN": "6", "genetiker|NOUN": "6", "sextionde|NUM": "6", "timmerstock|NOUN": "6", "bjälke|NOUN": "6", "excellens|NOUN": "6", "läsesal|NOUN": "6", "profylax|NOUN": "6", "koordinator|NOUN": "6", "poängställning|NOUN": "6", "docka|VERB": "6", "fjärran|NOUN": "6", "territorial|ADJ": "6", "grafiker|NOUN": "6", "undertröja|NOUN": "6", "anfallsspelare|NOUN": "6", "blotta|NOUN": "6", "förfrågan|NOUN": "6", "raffinera|VERB": "6", "specificitet|NOUN": "6", "begeistring|NOUN": "6", "bergskam|NOUN": "6", "okultiverad|ADJ": "6", "skrynkla|NOUN": "6", "statistiker|NOUN": "6", "syra|VERB": "6", "vinäger|NOUN": "6", "upphetsa|VERB": "6", "författningsenlig|ADJ": "6", "kalsong|NOUN": "6", "klagan|NOUN": "6", "kvitt|NOUN": "6", "planta|VERB": "6", "toppen|ADJ": "6", "tvåsidig|ADJ": "6"}